library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ALPR_constants is

  constant c_TEMPLATE_MASK : std_logic_vector(3999 downto 0) := x"0x3fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc00003fffffffffffffffffffc0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

end ALPR_constants;
