library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Package_Fixed.all;

package Package_Constant is

------------------------------------ 16 bits (8.8) -----------------------------------
--   constant c_Gaussian_Kernel_3 : fixed_vector(8 downto 0) := (
--     0=> x"0013", 1=> x"0020", 2=> x"0013",
--     3=> x"0020", 4=> x"0034", 5=> x"0020",
--     6=> x"0013", 7=> x"0020", 8=> x"0013"
--   );
--
--   constant c_Gaussian_Kernel_5 : fixed_vector(24 downto 0) := (
--     0=> x"0001",  1=> x"0003",  2=> x"0006",  3=> x"0003",  4=> x"0001",
--     5=> x"0003",  6=> x"000f",  7=> x"0019",  8=> x"000f",  9=> x"0003",
--     10=> x"0006", 11=> x"0019", 12=> x"0029", 13=> x"0019", 14=> x"0006",
--     15=> x"0003", 16=> x"000f", 17=> x"0019", 18=> x"000f", 19=> x"0003",
--     20=> x"0001", 21=> x"0003", 22=> x"0006", 23=> x"0003", 24=> x"0001"
--   );
--
--   constant c_Gaussian_Kernel_7 : fixed_vector(48 downto 0) := (
--     0=> x"0000",  1=> x"0000", 2=> x"0000",  3=> x"0000",   4=> x"0000",  5=> x"0000",  6=> x"0000",
--     7=> x"0000",  8=> x"0001", 9=> x"0003",  10=> x"0006",  11=> x"0003", 12=> x"0001", 13=> x"0000",
--     14=> x"0000", 15=> x"0003", 16=> x"000f", 17=> x"0019", 18=> x"000f", 19=> x"0003", 20=> x"0000",
--     21=> x"0000", 22=> x"0006", 23=> x"0019", 24=> x"0029", 25=> x"0019", 26=> x"0006", 27=> x"0000",
--     28=> x"0000", 29=> x"0003", 30=> x"000f", 31=> x"0019", 32=> x"000f", 33=> x"0003", 34=> x"0000",
--     35=> x"0000", 36=> x"0001", 37=> x"0003", 38=> x"0006", 39=> x"0003", 40=> x"0001", 41=> x"0000",
--     42=> x"0000", 43=> x"0000", 44=> x"0000", 45=> x"0000", 46=> x"0000", 47=> x"0000", 48=> x"0000"
--   );
-- ------------------------------------ 18 bits (10.8)  -----------------------------------
--   -- constant c_Gaussian_Kernel_3 : fixed_vector(8 downto 0) := (
--   --   0=>"0000000000000010011", 1=>"0000000000000100000", 2=>"0000000000000010011",
--   --   3=>"0000000000000100000", 4=>"0000000000000110100", 5=>"0000000000000100000",
--   --   6=>"0000000000000010011", 7=>"0000000000000100000", 8=>"0000000000000010011"
--   -- );
--   -- -- 19 bits (11.8)
--   -- constant c_Gaussian_Kernel_5 : fixed_vector(24 downto 0) := (
--   -- 0=>"0000000000000000001",  1=>"0000000000000000011",  2=>"0000000000000000110",  3=>"0000000000000000011",  4=>"0000000000000000001",
--   -- 5=>"0000000000000000011",  6=>"0000000000000001111",  7=>"0000000000000011001",  8=>"0000000000000001111",  9=>"0000000000000000011",
--   -- 10=>"0000000000000000110", 11=>"0000000000000011001", 12=>"0000000000000101001", 13=>"0000000000000011001", 14=>"0000000000000000110",
--   -- 15=>"0000000000000000011", 16=>"0000000000000001111", 17=>"0000000000000011001", 18=>"0000000000000001111", 19=>"0000000000000000011",
--   -- 20=>"0000000000000000001", 21=>"0000000000000000011", 22=>"0000000000000000110", 23=>"0000000000000000011", 24=>"0000000000000000001"
--   -- );
--   --
--   -- constant c_Gaussian_Kernel_7 : fixed_vector(48 downto 0) := (
--   -- 0 =>"0000000000000000000",  1=>"0000000000000000000",  2=>"0000000000000000000",   3=>"0000000000000000000",  4=>"0000000000000000000",  5=>"0000000000000000000",  6=>"0000000000000000000",
--   -- 7=>"0000000000000000000",   8 =>"0000000000000000001",  9=>"0000000000000000011", 10=>"0000000000000000110", 11=>"0000000000000000011", 12=>"0000000000000000001", 13=>"0000000000000000000",
--   -- 14=>"0000000000000000000",  15=>"0000000000000000011", 16=>"0000000000000001111", 17=>"0000000000000011001", 18=>"0000000000000001111", 19=>"0000000000000000011", 20=>"0000000000000000000",
--   -- 21=>"0000000000000000000",  22=>"0000000000000000110", 23=>"0000000000000011001", 24=>"0000000000000101001", 25=>"0000000000000011001", 26=>"0000000000000000110", 27=>"0000000000000000000",
--   -- 28=>"0000000000000000000",  29=>"0000000000000000011", 30=>"0000000000000001111", 31=>"0000000000000011001",  32=>"0000000000000001111", 33=>"0000000000000000011", 34=>"0000000000000000000",
--   -- 35=>"0000000000000000000",  36=>"0000000000000000001", 37=>"0000000000000000011", 38=>"0000000000000000110",  39=>"0000000000000000011", 40=>"0000000000000000001", 41=>"0000000000000000000",
--   -- 42=>"0000000000000000000",  43=>"0000000000000000000", 44=>"0000000000000000000", 45=>"0000000000000000000",  46=>"0000000000000000000", 47=>"0000000000000000000", 48=>"0000000000000000000"
--   -- );
-- ------------------------------------ 12 bits (8.4) -----------------------------------
--   -- constant c_Gaussian_Kernel_3 : fixed_vector(8 downto 0) := (
--   --   0=> x"001", 1=> x"002", 2=> x"001",
--   --   3=> x"002", 4=> x"003", 5=> x"002",
--   --   6=> x"001", 7=> x"002", 8=> x"001"
--   -- );
--   --
--   -- constant c_Gaussian_Kernel_5 : fixed_vector(24 downto 0) := (
--   --   0=>   x"000", 1=>   x"000", 2=>   x"000", 3=>   x"000", 4=>   x"000",
--   --   5=>   x"000", 6=>   x"001", 7=>   x"002", 8=>   x"001", 9=>   x"000",
--   --   10=>  x"000", 11=>  x"002", 12=>  x"003", 13=>  x"002", 14=>  x"000",
--   --   15=>  x"000", 16=>  x"001", 17=>  x"002", 18=>  x"001", 19=>  x"000",
--   --   20=>  x"000", 21=>  x"000", 22=>  x"000", 23=>  x"000", 24=>  x"000"
--   -- );
--   --
--   -- constant c_Gaussian_Kernel_7 : fixed_vector(48 downto 0) := (
--   --   0=>   x"000", 1=>   x"000", 2=>   x"000", 3=>   x"000", 4=>   x"000", 5=>   x"000", 6=>   x"000",
--   --   7=>   x"000", 8=>   x"000", 9=>   x"000", 10=>  x"000", 11=>  x"000", 12=>  x"000", 13=>  x"000",
--   --   14=>  x"000", 15=>  x"000", 16=>  x"001", 17=>  x"002", 18=>  x"001", 19=>  x"000", 20=>  x"000",
--   --   21=>  x"000", 22=>  x"000", 23=>  x"002", 24=>  x"003", 25=>  x"002", 26=>  x"000", 27=>  x"000",
--   --   28=>  x"000", 29=>  x"000", 30=>  x"001", 31=>  x"002", 32=>  x"001", 33=>  x"000", 34=>  x"000",
--   --   35=>  x"000", 36=>  x"000", 37=>  x"000", 38=>  x"000", 39=>  x"000", 40=>  x"000", 41=>  x"000",
--   --   42=>  x"000", 43=>  x"000", 44=>  x"000", 45=>  x"000", 46=>  x"000", 47=>  x"000", 48=>  x"000"
--   -- );
--
-- -------------------------------------- LUT constants ---------------------------
-- -- 3x3
-- constant c_Gaussian_Lut_3_W0: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0013",	2 => x"0026",	3 => x"0039",
-- 4 => x"004c",	5 => x"005f",	6 => x"0072",	7 => x"0085",
-- 8 => x"0098",	9 => x"00ab",	10 => x"00be",	11 => x"00d1",
-- 12 => x"00e4",	13 => x"00f7",	14 => x"010a",	15 => x"011d",
-- 16 => x"0130",	17 => x"0143",	18 => x"0156",	19 => x"0169",
-- 20 => x"017c",	21 => x"018f",	22 => x"01a2",	23 => x"01b5",
-- 24 => x"01c8",	25 => x"01db",	26 => x"01ee",	27 => x"0201",
-- 28 => x"0214",	29 => x"0227",	30 => x"023a",	31 => x"024d",
-- 32 => x"0260",	33 => x"0273",	34 => x"0286",	35 => x"0299",
-- 36 => x"02ac",	37 => x"02bf",	38 => x"02d2",	39 => x"02e5",
-- 40 => x"02f8",	41 => x"030b",	42 => x"031e",	43 => x"0331",
-- 44 => x"0344",	45 => x"0357",	46 => x"036a",	47 => x"037d",
-- 48 => x"0390",	49 => x"03a3",	50 => x"03b6",	51 => x"03c9",
-- 52 => x"03dc",	53 => x"03ef",	54 => x"0402",	55 => x"0415",
-- 56 => x"0428",	57 => x"043b",	58 => x"044e",	59 => x"0461",
-- 60 => x"0474",	61 => x"0487",	62 => x"049a",	63 => x"04ad",
-- 64 => x"04c0",	65 => x"04d3",	66 => x"04e6",	67 => x"04f9",
-- 68 => x"050c",	69 => x"051f",	70 => x"0532",	71 => x"0545",
-- 72 => x"0558",	73 => x"056b",	74 => x"057e",	75 => x"0591",
-- 76 => x"05a4",	77 => x"05b7",	78 => x"05ca",	79 => x"05dd",
-- 80 => x"05f0",	81 => x"0603",	82 => x"0616",	83 => x"0629",
-- 84 => x"063c",	85 => x"064f",	86 => x"0662",	87 => x"0675",
-- 88 => x"0688",	89 => x"069b",	90 => x"06ae",	91 => x"06c1",
-- 92 => x"06d4",	93 => x"06e7",	94 => x"06fa",	95 => x"070d",
-- 96 => x"0720",	97 => x"0733",	98 => x"0746",	99 => x"0759",
-- 100 => x"076c",	101 => x"077f",	102 => x"0792",	103 => x"07a5",
-- 104 => x"07b8",	105 => x"07cb",	106 => x"07de",	107 => x"07f1",
-- 108 => x"0804",	109 => x"0817",	110 => x"082a",	111 => x"083d",
-- 112 => x"0850",	113 => x"0863",	114 => x"0876",	115 => x"0889",
-- 116 => x"089c",	117 => x"08af",	118 => x"08c2",	119 => x"08d5",
-- 120 => x"08e8",	121 => x"08fb",	122 => x"090e",	123 => x"0921",
-- 124 => x"0934",	125 => x"0947",	126 => x"095a",	127 => x"096d",
-- 128 => x"0980",	129 => x"0993",	130 => x"09a6",	131 => x"09b9",
-- 132 => x"09cc",	133 => x"09df",	134 => x"09f2",	135 => x"0a05",
-- 136 => x"0a18",	137 => x"0a2b",	138 => x"0a3e",	139 => x"0a51",
-- 140 => x"0a64",	141 => x"0a77",	142 => x"0a8a",	143 => x"0a9d",
-- 144 => x"0ab0",	145 => x"0ac3",	146 => x"0ad6",	147 => x"0ae9",
-- 148 => x"0afc",	149 => x"0b0f",	150 => x"0b22",	151 => x"0b35",
-- 152 => x"0b48",	153 => x"0b5b",	154 => x"0b6e",	155 => x"0b81",
-- 156 => x"0b94",	157 => x"0ba7",	158 => x"0bba",	159 => x"0bcd",
-- 160 => x"0be0",	161 => x"0bf3",	162 => x"0c06",	163 => x"0c19",
-- 164 => x"0c2c",	165 => x"0c3f",	166 => x"0c52",	167 => x"0c65",
-- 168 => x"0c78",	169 => x"0c8b",	170 => x"0c9e",	171 => x"0cb1",
-- 172 => x"0cc4",	173 => x"0cd7",	174 => x"0cea",	175 => x"0cfd",
-- 176 => x"0d10",	177 => x"0d23",	178 => x"0d36",	179 => x"0d49",
-- 180 => x"0d5c",	181 => x"0d6f",	182 => x"0d82",	183 => x"0d95",
-- 184 => x"0da8",	185 => x"0dbb",	186 => x"0dce",	187 => x"0de1",
-- 188 => x"0df4",	189 => x"0e07",	190 => x"0e1a",	191 => x"0e2d",
-- 192 => x"0e40",	193 => x"0e53",	194 => x"0e66",	195 => x"0e79",
-- 196 => x"0e8c",	197 => x"0e9f",	198 => x"0eb2",	199 => x"0ec5",
-- 200 => x"0ed8",	201 => x"0eeb",	202 => x"0efe",	203 => x"0f11",
-- 204 => x"0f24",	205 => x"0f37",	206 => x"0f4a",	207 => x"0f5d",
-- 208 => x"0f70",	209 => x"0f83",	210 => x"0f96",	211 => x"0fa9",
-- 212 => x"0fbc",	213 => x"0fcf",	214 => x"0fe2",	215 => x"0ff5",
-- 216 => x"1008",	217 => x"101b",	218 => x"102e",	219 => x"1041",
-- 220 => x"1054",	221 => x"1067",	222 => x"107a",	223 => x"108d",
-- 224 => x"10a0",	225 => x"10b3",	226 => x"10c6",	227 => x"10d9",
-- 228 => x"10ec",	229 => x"10ff",	230 => x"1112",	231 => x"1125",
-- 232 => x"1138",	233 => x"114b",	234 => x"115e",	235 => x"1171",
-- 236 => x"1184",	237 => x"1197",	238 => x"11aa",	239 => x"11bd",
-- 240 => x"11d0",	241 => x"11e3",	242 => x"11f6",	243 => x"1209",
-- 244 => x"121c",	245 => x"122f",	246 => x"1242",	247 => x"1255",
-- 248 => x"1268",	249 => x"127b",	250 => x"128e",	251 => x"12a1",
-- 252 => x"12b4",	253 => x"12c7",	254 => x"12da",	255 => x"12ed");
--
-- constant c_Gaussian_Lut_3_W1: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0020",	2 => x"0040",	3 => x"0060",
-- 4 => x"0080",	5 => x"00a0",	6 => x"00c0",	7 => x"00e0",
-- 8 => x"0100",	9 => x"0120",	10 => x"0140",	11 => x"0160",
-- 12 => x"0180",	13 => x"01a0",	14 => x"01c0",	15 => x"01e0",
-- 16 => x"0200",	17 => x"0220",	18 => x"0240",	19 => x"0260",
-- 20 => x"0280",	21 => x"02a0",	22 => x"02c0",	23 => x"02e0",
-- 24 => x"0300",	25 => x"0320",	26 => x"0340",	27 => x"0360",
-- 28 => x"0380",	29 => x"03a0",	30 => x"03c0",	31 => x"03e0",
-- 32 => x"0400",	33 => x"0420",	34 => x"0440",	35 => x"0460",
-- 36 => x"0480",	37 => x"04a0",	38 => x"04c0",	39 => x"04e0",
-- 40 => x"0500",	41 => x"0520",	42 => x"0540",	43 => x"0560",
-- 44 => x"0580",	45 => x"05a0",	46 => x"05c0",	47 => x"05e0",
-- 48 => x"0600",	49 => x"0620",	50 => x"0640",	51 => x"0660",
-- 52 => x"0680",	53 => x"06a0",	54 => x"06c0",	55 => x"06e0",
-- 56 => x"0700",	57 => x"0720",	58 => x"0740",	59 => x"0760",
-- 60 => x"0780",	61 => x"07a0",	62 => x"07c0",	63 => x"07e0",
-- 64 => x"0800",	65 => x"0820",	66 => x"0840",	67 => x"0860",
-- 68 => x"0880",	69 => x"08a0",	70 => x"08c0",	71 => x"08e0",
-- 72 => x"0900",	73 => x"0920",	74 => x"0940",	75 => x"0960",
-- 76 => x"0980",	77 => x"09a0",	78 => x"09c0",	79 => x"09e0",
-- 80 => x"0a00",	81 => x"0a20",	82 => x"0a40",	83 => x"0a60",
-- 84 => x"0a80",	85 => x"0aa0",	86 => x"0ac0",	87 => x"0ae0",
-- 88 => x"0b00",	89 => x"0b20",	90 => x"0b40",	91 => x"0b60",
-- 92 => x"0b80",	93 => x"0ba0",	94 => x"0bc0",	95 => x"0be0",
-- 96 => x"0c00",	97 => x"0c20",	98 => x"0c40",	99 => x"0c60",
-- 100 => x"0c80",	101 => x"0ca0",	102 => x"0cc0",	103 => x"0ce0",
-- 104 => x"0d00",	105 => x"0d20",	106 => x"0d40",	107 => x"0d60",
-- 108 => x"0d80",	109 => x"0da0",	110 => x"0dc0",	111 => x"0de0",
-- 112 => x"0e00",	113 => x"0e20",	114 => x"0e40",	115 => x"0e60",
-- 116 => x"0e80",	117 => x"0ea0",	118 => x"0ec0",	119 => x"0ee0",
-- 120 => x"0f00",	121 => x"0f20",	122 => x"0f40",	123 => x"0f60",
-- 124 => x"0f80",	125 => x"0fa0",	126 => x"0fc0",	127 => x"0fe0",
-- 128 => x"1000",	129 => x"1020",	130 => x"1040",	131 => x"1060",
-- 132 => x"1080",	133 => x"10a0",	134 => x"10c0",	135 => x"10e0",
-- 136 => x"1100",	137 => x"1120",	138 => x"1140",	139 => x"1160",
-- 140 => x"1180",	141 => x"11a0",	142 => x"11c0",	143 => x"11e0",
-- 144 => x"1200",	145 => x"1220",	146 => x"1240",	147 => x"1260",
-- 148 => x"1280",	149 => x"12a0",	150 => x"12c0",	151 => x"12e0",
-- 152 => x"1300",	153 => x"1320",	154 => x"1340",	155 => x"1360",
-- 156 => x"1380",	157 => x"13a0",	158 => x"13c0",	159 => x"13e0",
-- 160 => x"1400",	161 => x"1420",	162 => x"1440",	163 => x"1460",
-- 164 => x"1480",	165 => x"14a0",	166 => x"14c0",	167 => x"14e0",
-- 168 => x"1500",	169 => x"1520",	170 => x"1540",	171 => x"1560",
-- 172 => x"1580",	173 => x"15a0",	174 => x"15c0",	175 => x"15e0",
-- 176 => x"1600",	177 => x"1620",	178 => x"1640",	179 => x"1660",
-- 180 => x"1680",	181 => x"16a0",	182 => x"16c0",	183 => x"16e0",
-- 184 => x"1700",	185 => x"1720",	186 => x"1740",	187 => x"1760",
-- 188 => x"1780",	189 => x"17a0",	190 => x"17c0",	191 => x"17e0",
-- 192 => x"1800",	193 => x"1820",	194 => x"1840",	195 => x"1860",
-- 196 => x"1880",	197 => x"18a0",	198 => x"18c0",	199 => x"18e0",
-- 200 => x"1900",	201 => x"1920",	202 => x"1940",	203 => x"1960",
-- 204 => x"1980",	205 => x"19a0",	206 => x"19c0",	207 => x"19e0",
-- 208 => x"1a00",	209 => x"1a20",	210 => x"1a40",	211 => x"1a60",
-- 212 => x"1a80",	213 => x"1aa0",	214 => x"1ac0",	215 => x"1ae0",
-- 216 => x"1b00",	217 => x"1b20",	218 => x"1b40",	219 => x"1b60",
-- 220 => x"1b80",	221 => x"1ba0",	222 => x"1bc0",	223 => x"1be0",
-- 224 => x"1c00",	225 => x"1c20",	226 => x"1c40",	227 => x"1c60",
-- 228 => x"1c80",	229 => x"1ca0",	230 => x"1cc0",	231 => x"1ce0",
-- 232 => x"1d00",	233 => x"1d20",	234 => x"1d40",	235 => x"1d60",
-- 236 => x"1d80",	237 => x"1da0",	238 => x"1dc0",	239 => x"1de0",
-- 240 => x"1e00",	241 => x"1e20",	242 => x"1e40",	243 => x"1e60",
-- 244 => x"1e80",	245 => x"1ea0",	246 => x"1ec0",	247 => x"1ee0",
-- 248 => x"1f00",	249 => x"1f20",	250 => x"1f40",	251 => x"1f60",
-- 252 => x"1f80",	253 => x"1fa0",	254 => x"1fc0",	255 => x"1fe0");
--
-- constant c_Gaussian_Lut_3_W2: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0034",	2 => x"0068",	3 => x"009c",
-- 4 => x"00d0",	5 => x"0104",	6 => x"0138",	7 => x"016c",
-- 8 => x"01a0",	9 => x"01d4",	10 => x"0208",	11 => x"023c",
-- 12 => x"0270",	13 => x"02a4",	14 => x"02d8",	15 => x"030c",
-- 16 => x"0340",	17 => x"0374",	18 => x"03a8",	19 => x"03dc",
-- 20 => x"0410",	21 => x"0444",	22 => x"0478",	23 => x"04ac",
-- 24 => x"04e0",	25 => x"0514",	26 => x"0548",	27 => x"057c",
-- 28 => x"05b0",	29 => x"05e4",	30 => x"0618",	31 => x"064c",
-- 32 => x"0680",	33 => x"06b4",	34 => x"06e8",	35 => x"071c",
-- 36 => x"0750",	37 => x"0784",	38 => x"07b8",	39 => x"07ec",
-- 40 => x"0820",	41 => x"0854",	42 => x"0888",	43 => x"08bc",
-- 44 => x"08f0",	45 => x"0924",	46 => x"0958",	47 => x"098c",
-- 48 => x"09c0",	49 => x"09f4",	50 => x"0a28",	51 => x"0a5c",
-- 52 => x"0a90",	53 => x"0ac4",	54 => x"0af8",	55 => x"0b2c",
-- 56 => x"0b60",	57 => x"0b94",	58 => x"0bc8",	59 => x"0bfc",
-- 60 => x"0c30",	61 => x"0c64",	62 => x"0c98",	63 => x"0ccc",
-- 64 => x"0d00",	65 => x"0d34",	66 => x"0d68",	67 => x"0d9c",
-- 68 => x"0dd0",	69 => x"0e04",	70 => x"0e38",	71 => x"0e6c",
-- 72 => x"0ea0",	73 => x"0ed4",	74 => x"0f08",	75 => x"0f3c",
-- 76 => x"0f70",	77 => x"0fa4",	78 => x"0fd8",	79 => x"100c",
-- 80 => x"1040",	81 => x"1074",	82 => x"10a8",	83 => x"10dc",
-- 84 => x"1110",	85 => x"1144",	86 => x"1178",	87 => x"11ac",
-- 88 => x"11e0",	89 => x"1214",	90 => x"1248",	91 => x"127c",
-- 92 => x"12b0",	93 => x"12e4",	94 => x"1318",	95 => x"134c",
-- 96 => x"1380",	97 => x"13b4",	98 => x"13e8",	99 => x"141c",
-- 100 => x"1450",	101 => x"1484",	102 => x"14b8",	103 => x"14ec",
-- 104 => x"1520",	105 => x"1554",	106 => x"1588",	107 => x"15bc",
-- 108 => x"15f0",	109 => x"1624",	110 => x"1658",	111 => x"168c",
-- 112 => x"16c0",	113 => x"16f4",	114 => x"1728",	115 => x"175c",
-- 116 => x"1790",	117 => x"17c4",	118 => x"17f8",	119 => x"182c",
-- 120 => x"1860",	121 => x"1894",	122 => x"18c8",	123 => x"18fc",
-- 124 => x"1930",	125 => x"1964",	126 => x"1998",	127 => x"19cc",
-- 128 => x"1a00",	129 => x"1a34",	130 => x"1a68",	131 => x"1a9c",
-- 132 => x"1ad0",	133 => x"1b04",	134 => x"1b38",	135 => x"1b6c",
-- 136 => x"1ba0",	137 => x"1bd4",	138 => x"1c08",	139 => x"1c3c",
-- 140 => x"1c70",	141 => x"1ca4",	142 => x"1cd8",	143 => x"1d0c",
-- 144 => x"1d40",	145 => x"1d74",	146 => x"1da8",	147 => x"1ddc",
-- 148 => x"1e10",	149 => x"1e44",	150 => x"1e78",	151 => x"1eac",
-- 152 => x"1ee0",	153 => x"1f14",	154 => x"1f48",	155 => x"1f7c",
-- 156 => x"1fb0",	157 => x"1fe4",	158 => x"2018",	159 => x"204c",
-- 160 => x"2080",	161 => x"20b4",	162 => x"20e8",	163 => x"211c",
-- 164 => x"2150",	165 => x"2184",	166 => x"21b8",	167 => x"21ec",
-- 168 => x"2220",	169 => x"2254",	170 => x"2288",	171 => x"22bc",
-- 172 => x"22f0",	173 => x"2324",	174 => x"2358",	175 => x"238c",
-- 176 => x"23c0",	177 => x"23f4",	178 => x"2428",	179 => x"245c",
-- 180 => x"2490",	181 => x"24c4",	182 => x"24f8",	183 => x"252c",
-- 184 => x"2560",	185 => x"2594",	186 => x"25c8",	187 => x"25fc",
-- 188 => x"2630",	189 => x"2664",	190 => x"2698",	191 => x"26cc",
-- 192 => x"2700",	193 => x"2734",	194 => x"2768",	195 => x"279c",
-- 196 => x"27d0",	197 => x"2804",	198 => x"2838",	199 => x"286c",
-- 200 => x"28a0",	201 => x"28d4",	202 => x"2908",	203 => x"293c",
-- 204 => x"2970",	205 => x"29a4",	206 => x"29d8",	207 => x"2a0c",
-- 208 => x"2a40",	209 => x"2a74",	210 => x"2aa8",	211 => x"2adc",
-- 212 => x"2b10",	213 => x"2b44",	214 => x"2b78",	215 => x"2bac",
-- 216 => x"2be0",	217 => x"2c14",	218 => x"2c48",	219 => x"2c7c",
-- 220 => x"2cb0",	221 => x"2ce4",	222 => x"2d18",	223 => x"2d4c",
-- 224 => x"2d80",	225 => x"2db4",	226 => x"2de8",	227 => x"2e1c",
-- 228 => x"2e50",	229 => x"2e84",	230 => x"2eb8",	231 => x"2eec",
-- 232 => x"2f20",	233 => x"2f54",	234 => x"2f88",	235 => x"2fbc",
-- 236 => x"2ff0",	237 => x"3024",	238 => x"3058",	239 => x"308c",
-- 240 => x"30c0",	241 => x"30f4",	242 => x"3128",	243 => x"315c",
-- 244 => x"3190",	245 => x"31c4",	246 => x"31f8",	247 => x"322c",
-- 248 => x"3260",	249 => x"3294",	250 => x"32c8",	251 => x"32fc",
-- 252 => x"3330",	253 => x"3364",	254 => x"3398",	255 => x"33cc");
--
-- --5x5
-- constant c_Gaussian_Lut_5_W0: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0001",	2 => x"0002",	3 => x"0003",	4 => x"0004",	5 => x"0005",
-- 6 => x"0006",	7 => x"0007",	8 => x"0008",	9 => x"0009",	10 => x"000a",	11 => x"000b",
-- 12 => x"000c",	13 => x"000d",	14 => x"000e",	15 => x"000f",	16 => x"0010",	17 => x"0011",
-- 18 => x"0012",	19 => x"0013",	20 => x"0014",	21 => x"0015",	22 => x"0016",	23 => x"0017",
-- 24 => x"0018",	25 => x"0019",	26 => x"001a",	27 => x"001b",	28 => x"001c",	29 => x"001d",
-- 30 => x"001e",	31 => x"001f",	32 => x"0020",	33 => x"0021",	34 => x"0022",	35 => x"0023",
-- 36 => x"0024",	37 => x"0025",	38 => x"0026",	39 => x"0027",	40 => x"0028",	41 => x"0029",
-- 42 => x"002a",	43 => x"002b",	44 => x"002c",	45 => x"002d",	46 => x"002e",	47 => x"002f",
-- 48 => x"0030",	49 => x"0031",	50 => x"0032",	51 => x"0033",	52 => x"0034",	53 => x"0035",
-- 54 => x"0036",	55 => x"0037",	56 => x"0038",	57 => x"0039",	58 => x"003a",	59 => x"003b",
-- 60 => x"003c",	61 => x"003d",	62 => x"003e",	63 => x"003f",	64 => x"0040",	65 => x"0041",
-- 66 => x"0042",	67 => x"0043",	68 => x"0044",	69 => x"0045",	70 => x"0046",	71 => x"0047",
-- 72 => x"0048",	73 => x"0049",	74 => x"004a",	75 => x"004b",	76 => x"004c",	77 => x"004d",
-- 78 => x"004e",	79 => x"004f",	80 => x"0050",	81 => x"0051",	82 => x"0052",	83 => x"0053",
-- 84 => x"0054",	85 => x"0055",	86 => x"0056",	87 => x"0057",	88 => x"0058",	89 => x"0059",
-- 90 => x"005a",	91 => x"005b",	92 => x"005c",	93 => x"005d",	94 => x"005e",	95 => x"005f",
-- 96 => x"0060",	97 => x"0061",	98 => x"0062",	99 => x"0063",	100 => x"0064",	101 => x"0065",
-- 102 => x"0066",	103 => x"0067",	104 => x"0068",	105 => x"0069",	106 => x"006a",	107 => x"006b",
-- 108 => x"006c",	109 => x"006d",	110 => x"006e",	111 => x"006f",	112 => x"0070",	113 => x"0071",
-- 114 => x"0072",	115 => x"0073",	116 => x"0074",	117 => x"0075",	118 => x"0076",	119 => x"0077",
-- 120 => x"0078",	121 => x"0079",	122 => x"007a",	123 => x"007b",	124 => x"007c",	125 => x"007d",
-- 126 => x"007e",	127 => x"007f",	128 => x"0080",	129 => x"0081",	130 => x"0082",	131 => x"0083",
-- 132 => x"0084",	133 => x"0085",	134 => x"0086",	135 => x"0087",	136 => x"0088",	137 => x"0089",
-- 138 => x"008a",	139 => x"008b",	140 => x"008c",	141 => x"008d",	142 => x"008e",	143 => x"008f",
-- 144 => x"0090",	145 => x"0091",	146 => x"0092",	147 => x"0093",	148 => x"0094",	149 => x"0095",
-- 150 => x"0096",	151 => x"0097",	152 => x"0098",	153 => x"0099",	154 => x"009a",	155 => x"009b",
-- 156 => x"009c",	157 => x"009d",	158 => x"009e",	159 => x"009f",	160 => x"00a0",	161 => x"00a1",
-- 162 => x"00a2",	163 => x"00a3",	164 => x"00a4",	165 => x"00a5",	166 => x"00a6",	167 => x"00a7",
-- 168 => x"00a8",	169 => x"00a9",	170 => x"00aa",	171 => x"00ab",	172 => x"00ac",	173 => x"00ad",
-- 174 => x"00ae",	175 => x"00af",	176 => x"00b0",	177 => x"00b1",	178 => x"00b2",	179 => x"00b3",
-- 180 => x"00b4",	181 => x"00b5",	182 => x"00b6",	183 => x"00b7",	184 => x"00b8",	185 => x"00b9",
-- 186 => x"00ba",	187 => x"00bb",	188 => x"00bc",	189 => x"00bd",	190 => x"00be",	191 => x"00bf",
-- 192 => x"00c0",	193 => x"00c1",	194 => x"00c2",	195 => x"00c3",	196 => x"00c4",	197 => x"00c5",
-- 198 => x"00c6",	199 => x"00c7",	200 => x"00c8",	201 => x"00c9",	202 => x"00ca",	203 => x"00cb",
-- 204 => x"00cc",	205 => x"00cd",	206 => x"00ce",	207 => x"00cf",	208 => x"00d0",	209 => x"00d1",
-- 210 => x"00d2",	211 => x"00d3",	212 => x"00d4",	213 => x"00d5",	214 => x"00d6",	215 => x"00d7",
-- 216 => x"00d8",	217 => x"00d9",	218 => x"00da",	219 => x"00db",	220 => x"00dc",	221 => x"00dd",
-- 222 => x"00de",	223 => x"00df",	224 => x"00e0",	225 => x"00e1",	226 => x"00e2",	227 => x"00e3",
-- 228 => x"00e4",	229 => x"00e5",	230 => x"00e6",	231 => x"00e7",	232 => x"00e8",	233 => x"00e9",
-- 234 => x"00ea",	235 => x"00eb",	236 => x"00ec",	237 => x"00ed",	238 => x"00ee",	239 => x"00ef",
-- 240 => x"00f0",	241 => x"00f1",	242 => x"00f2",	243 => x"00f3",	244 => x"00f4",	245 => x"00f5",
-- 246 => x"00f6",	247 => x"00f7",	248 => x"00f8",	249 => x"00f9",	250 => x"00fa",	251 => x"00fb",
-- 252 => x"00fc",	253 => x"00fd",	254 => x"00fe",	255 => x"00ff");
--
-- constant c_Gaussian_Lut_5_W1: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0003",	2 => x"0006",	3 => x"0009",	4 => x"000c",	5 => x"000f",
-- 6 => x"0012",	7 => x"0015",	8 => x"0018",	9 => x"001b",	10 => x"001e",	11 => x"0021",
-- 12 => x"0024",	13 => x"0027",	14 => x"002a",	15 => x"002d",	16 => x"0030",	17 => x"0033",
-- 18 => x"0036",	19 => x"0039",	20 => x"003c",	21 => x"003f",	22 => x"0042",	23 => x"0045",
-- 24 => x"0048",	25 => x"004b",	26 => x"004e",	27 => x"0051",	28 => x"0054",	29 => x"0057",
-- 30 => x"005a",	31 => x"005d",	32 => x"0060",	33 => x"0063",	34 => x"0066",	35 => x"0069",
-- 36 => x"006c",	37 => x"006f",	38 => x"0072",	39 => x"0075",	40 => x"0078",	41 => x"007b",
-- 42 => x"007e",	43 => x"0081",	44 => x"0084",	45 => x"0087",	46 => x"008a",	47 => x"008d",
-- 48 => x"0090",	49 => x"0093",	50 => x"0096",	51 => x"0099",	52 => x"009c",	53 => x"009f",
-- 54 => x"00a2",	55 => x"00a5",	56 => x"00a8",	57 => x"00ab",	58 => x"00ae",	59 => x"00b1",
-- 60 => x"00b4",	61 => x"00b7",	62 => x"00ba",	63 => x"00bd",	64 => x"00c0",	65 => x"00c3",
-- 66 => x"00c6",	67 => x"00c9",	68 => x"00cc",	69 => x"00cf",	70 => x"00d2",	71 => x"00d5",
-- 72 => x"00d8",	73 => x"00db",	74 => x"00de",	75 => x"00e1",	76 => x"00e4",	77 => x"00e7",
-- 78 => x"00ea",	79 => x"00ed",	80 => x"00f0",	81 => x"00f3",	82 => x"00f6",	83 => x"00f9",
-- 84 => x"00fc",	85 => x"00ff",	86 => x"0102",	87 => x"0105",	88 => x"0108",	89 => x"010b",
-- 90 => x"010e",	91 => x"0111",	92 => x"0114",	93 => x"0117",	94 => x"011a",	95 => x"011d",
-- 96 => x"0120",	97 => x"0123",	98 => x"0126",	99 => x"0129",	100 => x"012c",	101 => x"012f",
-- 102 => x"0132",	103 => x"0135",	104 => x"0138",	105 => x"013b",	106 => x"013e",	107 => x"0141",
-- 108 => x"0144",	109 => x"0147",	110 => x"014a",	111 => x"014d",	112 => x"0150",	113 => x"0153",
-- 114 => x"0156",	115 => x"0159",	116 => x"015c",	117 => x"015f",	118 => x"0162",	119 => x"0165",
-- 120 => x"0168",	121 => x"016b",	122 => x"016e",	123 => x"0171",	124 => x"0174",	125 => x"0177",
-- 126 => x"017a",	127 => x"017d",	128 => x"0180",	129 => x"0183",	130 => x"0186",	131 => x"0189",
-- 132 => x"018c",	133 => x"018f",	134 => x"0192",	135 => x"0195",	136 => x"0198",	137 => x"019b",
-- 138 => x"019e",	139 => x"01a1",	140 => x"01a4",	141 => x"01a7",	142 => x"01aa",	143 => x"01ad",
-- 144 => x"01b0",	145 => x"01b3",	146 => x"01b6",	147 => x"01b9",	148 => x"01bc",	149 => x"01bf",
-- 150 => x"01c2",	151 => x"01c5",	152 => x"01c8",	153 => x"01cb",	154 => x"01ce",	155 => x"01d1",
-- 156 => x"01d4",	157 => x"01d7",	158 => x"01da",	159 => x"01dd",	160 => x"01e0",	161 => x"01e3",
-- 162 => x"01e6",	163 => x"01e9",	164 => x"01ec",	165 => x"01ef",	166 => x"01f2",	167 => x"01f5",
-- 168 => x"01f8",	169 => x"01fb",	170 => x"01fe",	171 => x"0201",	172 => x"0204",	173 => x"0207",
-- 174 => x"020a",	175 => x"020d",	176 => x"0210",	177 => x"0213",	178 => x"0216",	179 => x"0219",
-- 180 => x"021c",	181 => x"021f",	182 => x"0222",	183 => x"0225",	184 => x"0228",	185 => x"022b",
-- 186 => x"022e",	187 => x"0231",	188 => x"0234",	189 => x"0237",	190 => x"023a",	191 => x"023d",
-- 192 => x"0240",	193 => x"0243",	194 => x"0246",	195 => x"0249",	196 => x"024c",	197 => x"024f",
-- 198 => x"0252",	199 => x"0255",	200 => x"0258",	201 => x"025b",	202 => x"025e",	203 => x"0261",
-- 204 => x"0264",	205 => x"0267",	206 => x"026a",	207 => x"026d",	208 => x"0270",	209 => x"0273",
-- 210 => x"0276",	211 => x"0279",	212 => x"027c",	213 => x"027f",	214 => x"0282",	215 => x"0285",
-- 216 => x"0288",	217 => x"028b",	218 => x"028e",	219 => x"0291",	220 => x"0294",	221 => x"0297",
-- 222 => x"029a",	223 => x"029d",	224 => x"02a0",	225 => x"02a3",	226 => x"02a6",	227 => x"02a9",
-- 228 => x"02ac",	229 => x"02af",	230 => x"02b2",	231 => x"02b5",	232 => x"02b8",	233 => x"02bb",
-- 234 => x"02be",	235 => x"02c1",	236 => x"02c4",	237 => x"02c7",	238 => x"02ca",	239 => x"02cd",
-- 240 => x"02d0",	241 => x"02d3",	242 => x"02d6",	243 => x"02d9",	244 => x"02dc",	245 => x"02df",
-- 246 => x"02e2",	247 => x"02e5",	248 => x"02e8",	249 => x"02eb",	250 => x"02ee",	251 => x"02f1",
-- 252 => x"02f4",	253 => x"02f7",	254 => x"02fa",	255 => x"02fd");
--
-- constant c_Gaussian_Lut_5_W2: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0006",	2 => x"000c",	3 => x"0012",	4 => x"0018",	5 => x"001e",
-- 6 => x"0024",	7 => x"002a",	8 => x"0030",	9 => x"0036",	10 => x"003c",	11 => x"0042",
-- 12 => x"0048",	13 => x"004e",	14 => x"0054",	15 => x"005a",	16 => x"0060",	17 => x"0066",
-- 18 => x"006c",	19 => x"0072",	20 => x"0078",	21 => x"007e",	22 => x"0084",	23 => x"008a",
-- 24 => x"0090",	25 => x"0096",	26 => x"009c",	27 => x"00a2",	28 => x"00a8",	29 => x"00ae",
-- 30 => x"00b4",	31 => x"00ba",	32 => x"00c0",	33 => x"00c6",	34 => x"00cc",	35 => x"00d2",
-- 36 => x"00d8",	37 => x"00de",	38 => x"00e4",	39 => x"00ea",	40 => x"00f0",	41 => x"00f6",
-- 42 => x"00fc",	43 => x"0102",	44 => x"0108",	45 => x"010e",	46 => x"0114",	47 => x"011a",
-- 48 => x"0120",	49 => x"0126",	50 => x"012c",	51 => x"0132",	52 => x"0138",	53 => x"013e",
-- 54 => x"0144",	55 => x"014a",	56 => x"0150",	57 => x"0156",	58 => x"015c",	59 => x"0162",
-- 60 => x"0168",	61 => x"016e",	62 => x"0174",	63 => x"017a",	64 => x"0180",	65 => x"0186",
-- 66 => x"018c",	67 => x"0192",	68 => x"0198",	69 => x"019e",	70 => x"01a4",	71 => x"01aa",
-- 72 => x"01b0",	73 => x"01b6",	74 => x"01bc",	75 => x"01c2",	76 => x"01c8",	77 => x"01ce",
-- 78 => x"01d4",	79 => x"01da",	80 => x"01e0",	81 => x"01e6",	82 => x"01ec",	83 => x"01f2",
-- 84 => x"01f8",	85 => x"01fe",	86 => x"0204",	87 => x"020a",	88 => x"0210",	89 => x"0216",
-- 90 => x"021c",	91 => x"0222",	92 => x"0228",	93 => x"022e",	94 => x"0234",	95 => x"023a",
-- 96 => x"0240",	97 => x"0246",	98 => x"024c",	99 => x"0252",	100 => x"0258",	101 => x"025e",
-- 102 => x"0264",	103 => x"026a",	104 => x"0270",	105 => x"0276",	106 => x"027c",	107 => x"0282",
-- 108 => x"0288",	109 => x"028e",	110 => x"0294",	111 => x"029a",	112 => x"02a0",	113 => x"02a6",
-- 114 => x"02ac",	115 => x"02b2",	116 => x"02b8",	117 => x"02be",	118 => x"02c4",	119 => x"02ca",
-- 120 => x"02d0",	121 => x"02d6",	122 => x"02dc",	123 => x"02e2",	124 => x"02e8",	125 => x"02ee",
-- 126 => x"02f4",	127 => x"02fa",	128 => x"0300",	129 => x"0306",	130 => x"030c",	131 => x"0312",
-- 132 => x"0318",	133 => x"031e",	134 => x"0324",	135 => x"032a",	136 => x"0330",	137 => x"0336",
-- 138 => x"033c",	139 => x"0342",	140 => x"0348",	141 => x"034e",	142 => x"0354",	143 => x"035a",
-- 144 => x"0360",	145 => x"0366",	146 => x"036c",	147 => x"0372",	148 => x"0378",	149 => x"037e",
-- 150 => x"0384",	151 => x"038a",	152 => x"0390",	153 => x"0396",	154 => x"039c",	155 => x"03a2",
-- 156 => x"03a8",	157 => x"03ae",	158 => x"03b4",	159 => x"03ba",	160 => x"03c0",	161 => x"03c6",
-- 162 => x"03cc",	163 => x"03d2",	164 => x"03d8",	165 => x"03de",	166 => x"03e4",	167 => x"03ea",
-- 168 => x"03f0",	169 => x"03f6",	170 => x"03fc",	171 => x"0402",	172 => x"0408",	173 => x"040e",
-- 174 => x"0414",	175 => x"041a",	176 => x"0420",	177 => x"0426",	178 => x"042c",	179 => x"0432",
-- 180 => x"0438",	181 => x"043e",	182 => x"0444",	183 => x"044a",	184 => x"0450",	185 => x"0456",
-- 186 => x"045c",	187 => x"0462",	188 => x"0468",	189 => x"046e",	190 => x"0474",	191 => x"047a",
-- 192 => x"0480",	193 => x"0486",	194 => x"048c",	195 => x"0492",	196 => x"0498",	197 => x"049e",
-- 198 => x"04a4",	199 => x"04aa",	200 => x"04b0",	201 => x"04b6",	202 => x"04bc",	203 => x"04c2",
-- 204 => x"04c8",	205 => x"04ce",	206 => x"04d4",	207 => x"04da",	208 => x"04e0",	209 => x"04e6",
-- 210 => x"04ec",	211 => x"04f2",	212 => x"04f8",	213 => x"04fe",	214 => x"0504",	215 => x"050a",
-- 216 => x"0510",	217 => x"0516",	218 => x"051c",	219 => x"0522",	220 => x"0528",	221 => x"052e",
-- 222 => x"0534",	223 => x"053a",	224 => x"0540",	225 => x"0546",	226 => x"054c",	227 => x"0552",
-- 228 => x"0558",	229 => x"055e",	230 => x"0564",	231 => x"056a",	232 => x"0570",	233 => x"0576",
-- 234 => x"057c",	235 => x"0582",	236 => x"0588",	237 => x"058e",	238 => x"0594",	239 => x"059a",
-- 240 => x"05a0",	241 => x"05a6",	242 => x"05ac",	243 => x"05b2",	244 => x"05b8",	245 => x"05be",
-- 246 => x"05c4",	247 => x"05ca",	248 => x"05d0",	249 => x"05d6",	250 => x"05dc",	251 => x"05e2",
-- 252 => x"05e8",	253 => x"05ee",	254 => x"05f4",	255 => x"05fa");
--
-- constant c_Gaussian_Lut_5_W3: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"000f",	2 => x"001e",	3 => x"002d",	4 => x"003c",	5 => x"004b",
-- 6 => x"005a",	7 => x"0069",	8 => x"0078",	9 => x"0087",	10 => x"0096",	11 => x"00a5",
-- 12 => x"00b4",	13 => x"00c3",	14 => x"00d2",	15 => x"00e1",	16 => x"00f0",	17 => x"00ff",
-- 18 => x"010e",	19 => x"011d",	20 => x"012c",	21 => x"013b",	22 => x"014a",	23 => x"0159",
-- 24 => x"0168",	25 => x"0177",	26 => x"0186",	27 => x"0195",	28 => x"01a4",	29 => x"01b3",
-- 30 => x"01c2",	31 => x"01d1",	32 => x"01e0",	33 => x"01ef",	34 => x"01fe",	35 => x"020d",
-- 36 => x"021c",	37 => x"022b",	38 => x"023a",	39 => x"0249",	40 => x"0258",	41 => x"0267",
-- 42 => x"0276",	43 => x"0285",	44 => x"0294",	45 => x"02a3",	46 => x"02b2",	47 => x"02c1",
-- 48 => x"02d0",	49 => x"02df",	50 => x"02ee",	51 => x"02fd",	52 => x"030c",	53 => x"031b",
-- 54 => x"032a",	55 => x"0339",	56 => x"0348",	57 => x"0357",	58 => x"0366",	59 => x"0375",
-- 60 => x"0384",	61 => x"0393",	62 => x"03a2",	63 => x"03b1",	64 => x"03c0",	65 => x"03cf",
-- 66 => x"03de",	67 => x"03ed",	68 => x"03fc",	69 => x"040b",	70 => x"041a",	71 => x"0429",
-- 72 => x"0438",	73 => x"0447",	74 => x"0456",	75 => x"0465",	76 => x"0474",	77 => x"0483",
-- 78 => x"0492",	79 => x"04a1",	80 => x"04b0",	81 => x"04bf",	82 => x"04ce",	83 => x"04dd",
-- 84 => x"04ec",	85 => x"04fb",	86 => x"050a",	87 => x"0519",	88 => x"0528",	89 => x"0537",
-- 90 => x"0546",	91 => x"0555",	92 => x"0564",	93 => x"0573",	94 => x"0582",	95 => x"0591",
-- 96 => x"05a0",	97 => x"05af",	98 => x"05be",	99 => x"05cd",	100 => x"05dc",	101 => x"05eb",
-- 102 => x"05fa",	103 => x"0609",	104 => x"0618",	105 => x"0627",	106 => x"0636",	107 => x"0645",
-- 108 => x"0654",	109 => x"0663",	110 => x"0672",	111 => x"0681",	112 => x"0690",	113 => x"069f",
-- 114 => x"06ae",	115 => x"06bd",	116 => x"06cc",	117 => x"06db",	118 => x"06ea",	119 => x"06f9",
-- 120 => x"0708",	121 => x"0717",	122 => x"0726",	123 => x"0735",	124 => x"0744",	125 => x"0753",
-- 126 => x"0762",	127 => x"0771",	128 => x"0780",	129 => x"078f",	130 => x"079e",	131 => x"07ad",
-- 132 => x"07bc",	133 => x"07cb",	134 => x"07da",	135 => x"07e9",	136 => x"07f8",	137 => x"0807",
-- 138 => x"0816",	139 => x"0825",	140 => x"0834",	141 => x"0843",	142 => x"0852",	143 => x"0861",
-- 144 => x"0870",	145 => x"087f",	146 => x"088e",	147 => x"089d",	148 => x"08ac",	149 => x"08bb",
-- 150 => x"08ca",	151 => x"08d9",	152 => x"08e8",	153 => x"08f7",	154 => x"0906",	155 => x"0915",
-- 156 => x"0924",	157 => x"0933",	158 => x"0942",	159 => x"0951",	160 => x"0960",	161 => x"096f",
-- 162 => x"097e",	163 => x"098d",	164 => x"099c",	165 => x"09ab",	166 => x"09ba",	167 => x"09c9",
-- 168 => x"09d8",	169 => x"09e7",	170 => x"09f6",	171 => x"0a05",	172 => x"0a14",	173 => x"0a23",
-- 174 => x"0a32",	175 => x"0a41",	176 => x"0a50",	177 => x"0a5f",	178 => x"0a6e",	179 => x"0a7d",
-- 180 => x"0a8c",	181 => x"0a9b",	182 => x"0aaa",	183 => x"0ab9",	184 => x"0ac8",	185 => x"0ad7",
-- 186 => x"0ae6",	187 => x"0af5",	188 => x"0b04",	189 => x"0b13",	190 => x"0b22",	191 => x"0b31",
-- 192 => x"0b40",	193 => x"0b4f",	194 => x"0b5e",	195 => x"0b6d",	196 => x"0b7c",	197 => x"0b8b",
-- 198 => x"0b9a",	199 => x"0ba9",	200 => x"0bb8",	201 => x"0bc7",	202 => x"0bd6",	203 => x"0be5",
-- 204 => x"0bf4",	205 => x"0c03",	206 => x"0c12",	207 => x"0c21",	208 => x"0c30",	209 => x"0c3f",
-- 210 => x"0c4e",	211 => x"0c5d",	212 => x"0c6c",	213 => x"0c7b",	214 => x"0c8a",	215 => x"0c99",
-- 216 => x"0ca8",	217 => x"0cb7",	218 => x"0cc6",	219 => x"0cd5",	220 => x"0ce4",	221 => x"0cf3",
-- 222 => x"0d02",	223 => x"0d11",	224 => x"0d20",	225 => x"0d2f",	226 => x"0d3e",	227 => x"0d4d",
-- 228 => x"0d5c",	229 => x"0d6b",	230 => x"0d7a",	231 => x"0d89",	232 => x"0d98",	233 => x"0da7",
-- 234 => x"0db6",	235 => x"0dc5",	236 => x"0dd4",	237 => x"0de3",	238 => x"0df2",	239 => x"0e01",
-- 240 => x"0e10",	241 => x"0e1f",	242 => x"0e2e",	243 => x"0e3d",	244 => x"0e4c",	245 => x"0e5b",
-- 246 => x"0e6a",	247 => x"0e79",	248 => x"0e88",	249 => x"0e97",	250 => x"0ea6",	251 => x"0eb5",
-- 252 => x"0ec4",	253 => x"0ed3",	254 => x"0ee2",	255 => x"0ef1");
--
-- constant c_Gaussian_Lut_5_W4: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0019",	2 => x"0032",	3 => x"004b",	4 => x"0064",	5 => x"007d",
-- 6 => x"0096",	7 => x"00af",	8 => x"00c8",	9 => x"00e1",	10 => x"00fa",	11 => x"0113",
-- 12 => x"012c",	13 => x"0145",	14 => x"015e",	15 => x"0177",	16 => x"0190",	17 => x"01a9",
-- 18 => x"01c2",	19 => x"01db",	20 => x"01f4",	21 => x"020d",	22 => x"0226",	23 => x"023f",
-- 24 => x"0258",	25 => x"0271",	26 => x"028a",	27 => x"02a3",	28 => x"02bc",	29 => x"02d5",
-- 30 => x"02ee",	31 => x"0307",	32 => x"0320",	33 => x"0339",	34 => x"0352",	35 => x"036b",
-- 36 => x"0384",	37 => x"039d",	38 => x"03b6",	39 => x"03cf",	40 => x"03e8",	41 => x"0401",
-- 42 => x"041a",	43 => x"0433",	44 => x"044c",	45 => x"0465",	46 => x"047e",	47 => x"0497",
-- 48 => x"04b0",	49 => x"04c9",	50 => x"04e2",	51 => x"04fb",	52 => x"0514",	53 => x"052d",
-- 54 => x"0546",	55 => x"055f",	56 => x"0578",	57 => x"0591",	58 => x"05aa",	59 => x"05c3",
-- 60 => x"05dc",	61 => x"05f5",	62 => x"060e",	63 => x"0627",	64 => x"0640",	65 => x"0659",
-- 66 => x"0672",	67 => x"068b",	68 => x"06a4",	69 => x"06bd",	70 => x"06d6",	71 => x"06ef",
-- 72 => x"0708",	73 => x"0721",	74 => x"073a",	75 => x"0753",	76 => x"076c",	77 => x"0785",
-- 78 => x"079e",	79 => x"07b7",	80 => x"07d0",	81 => x"07e9",	82 => x"0802",	83 => x"081b",
-- 84 => x"0834",	85 => x"084d",	86 => x"0866",	87 => x"087f",	88 => x"0898",	89 => x"08b1",
-- 90 => x"08ca",	91 => x"08e3",	92 => x"08fc",	93 => x"0915",	94 => x"092e",	95 => x"0947",
-- 96 => x"0960",	97 => x"0979",	98 => x"0992",	99 => x"09ab",	100 => x"09c4",	101 => x"09dd",
-- 102 => x"09f6",	103 => x"0a0f",	104 => x"0a28",	105 => x"0a41",	106 => x"0a5a",	107 => x"0a73",
-- 108 => x"0a8c",	109 => x"0aa5",	110 => x"0abe",	111 => x"0ad7",	112 => x"0af0",	113 => x"0b09",
-- 114 => x"0b22",	115 => x"0b3b",	116 => x"0b54",	117 => x"0b6d",	118 => x"0b86",	119 => x"0b9f",
-- 120 => x"0bb8",	121 => x"0bd1",	122 => x"0bea",	123 => x"0c03",	124 => x"0c1c",	125 => x"0c35",
-- 126 => x"0c4e",	127 => x"0c67",	128 => x"0c80",	129 => x"0c99",	130 => x"0cb2",	131 => x"0ccb",
-- 132 => x"0ce4",	133 => x"0cfd",	134 => x"0d16",	135 => x"0d2f",	136 => x"0d48",	137 => x"0d61",
-- 138 => x"0d7a",	139 => x"0d93",	140 => x"0dac",	141 => x"0dc5",	142 => x"0dde",	143 => x"0df7",
-- 144 => x"0e10",	145 => x"0e29",	146 => x"0e42",	147 => x"0e5b",	148 => x"0e74",	149 => x"0e8d",
-- 150 => x"0ea6",	151 => x"0ebf",	152 => x"0ed8",	153 => x"0ef1",	154 => x"0f0a",	155 => x"0f23",
-- 156 => x"0f3c",	157 => x"0f55",	158 => x"0f6e",	159 => x"0f87",	160 => x"0fa0",	161 => x"0fb9",
-- 162 => x"0fd2",	163 => x"0feb",	164 => x"1004",	165 => x"101d",	166 => x"1036",	167 => x"104f",
-- 168 => x"1068",	169 => x"1081",	170 => x"109a",	171 => x"10b3",	172 => x"10cc",	173 => x"10e5",
-- 174 => x"10fe",	175 => x"1117",	176 => x"1130",	177 => x"1149",	178 => x"1162",	179 => x"117b",
-- 180 => x"1194",	181 => x"11ad",	182 => x"11c6",	183 => x"11df",	184 => x"11f8",	185 => x"1211",
-- 186 => x"122a",	187 => x"1243",	188 => x"125c",	189 => x"1275",	190 => x"128e",	191 => x"12a7",
-- 192 => x"12c0",	193 => x"12d9",	194 => x"12f2",	195 => x"130b",	196 => x"1324",	197 => x"133d",
-- 198 => x"1356",	199 => x"136f",	200 => x"1388",	201 => x"13a1",	202 => x"13ba",	203 => x"13d3",
-- 204 => x"13ec",	205 => x"1405",	206 => x"141e",	207 => x"1437",	208 => x"1450",	209 => x"1469",
-- 210 => x"1482",	211 => x"149b",	212 => x"14b4",	213 => x"14cd",	214 => x"14e6",	215 => x"14ff",
-- 216 => x"1518",	217 => x"1531",	218 => x"154a",	219 => x"1563",	220 => x"157c",	221 => x"1595",
-- 222 => x"15ae",	223 => x"15c7",	224 => x"15e0",	225 => x"15f9",	226 => x"1612",	227 => x"162b",
-- 228 => x"1644",	229 => x"165d",	230 => x"1676",	231 => x"168f",	232 => x"16a8",	233 => x"16c1",
-- 234 => x"16da",	235 => x"16f3",	236 => x"170c",	237 => x"1725",	238 => x"173e",	239 => x"1757",
-- 240 => x"1770",	241 => x"1789",	242 => x"17a2",	243 => x"17bb",	244 => x"17d4",	245 => x"17ed",
-- 246 => x"1806",	247 => x"181f",	248 => x"1838",	249 => x"1851",	250 => x"186a",	251 => x"1883",
-- 252 => x"189c",	253 => x"18b5",	254 => x"18ce",	255 => x"18e7");
--
-- constant c_Gaussian_Lut_5_W5: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0029",	2 => x"0052",	3 => x"007b",	4 => x"00a4",	5 => x"00cd",
-- 6 => x"00f6",	7 => x"011f",	8 => x"0148",	9 => x"0171",	10 => x"019a",	11 => x"01c3",
-- 12 => x"01ec",	13 => x"0215",	14 => x"023e",	15 => x"0267",	16 => x"0290",	17 => x"02b9",
-- 18 => x"02e2",	19 => x"030b",	20 => x"0334",	21 => x"035d",	22 => x"0386",	23 => x"03af",
-- 24 => x"03d8",	25 => x"0401",	26 => x"042a",	27 => x"0453",	28 => x"047c",	29 => x"04a5",
-- 30 => x"04ce",	31 => x"04f7",	32 => x"0520",	33 => x"0549",	34 => x"0572",	35 => x"059b",
-- 36 => x"05c4",	37 => x"05ed",	38 => x"0616",	39 => x"063f",	40 => x"0668",	41 => x"0691",
-- 42 => x"06ba",	43 => x"06e3",	44 => x"070c",	45 => x"0735",	46 => x"075e",	47 => x"0787",
-- 48 => x"07b0",	49 => x"07d9",	50 => x"0802",	51 => x"082b",	52 => x"0854",	53 => x"087d",
-- 54 => x"08a6",	55 => x"08cf",	56 => x"08f8",	57 => x"0921",	58 => x"094a",	59 => x"0973",
-- 60 => x"099c",	61 => x"09c5",	62 => x"09ee",	63 => x"0a17",	64 => x"0a40",	65 => x"0a69",
-- 66 => x"0a92",	67 => x"0abb",	68 => x"0ae4",	69 => x"0b0d",	70 => x"0b36",	71 => x"0b5f",
-- 72 => x"0b88",	73 => x"0bb1",	74 => x"0bda",	75 => x"0c03",	76 => x"0c2c",	77 => x"0c55",
-- 78 => x"0c7e",	79 => x"0ca7",	80 => x"0cd0",	81 => x"0cf9",	82 => x"0d22",	83 => x"0d4b",
-- 84 => x"0d74",	85 => x"0d9d",	86 => x"0dc6",	87 => x"0def",	88 => x"0e18",	89 => x"0e41",
-- 90 => x"0e6a",	91 => x"0e93",	92 => x"0ebc",	93 => x"0ee5",	94 => x"0f0e",	95 => x"0f37",
-- 96 => x"0f60",	97 => x"0f89",	98 => x"0fb2",	99 => x"0fdb",	100 => x"1004",	101 => x"102d",
-- 102 => x"1056",	103 => x"107f",	104 => x"10a8",	105 => x"10d1",	106 => x"10fa",	107 => x"1123",
-- 108 => x"114c",	109 => x"1175",	110 => x"119e",	111 => x"11c7",	112 => x"11f0",	113 => x"1219",
-- 114 => x"1242",	115 => x"126b",	116 => x"1294",	117 => x"12bd",	118 => x"12e6",	119 => x"130f",
-- 120 => x"1338",	121 => x"1361",	122 => x"138a",	123 => x"13b3",	124 => x"13dc",	125 => x"1405",
-- 126 => x"142e",	127 => x"1457",	128 => x"1480",	129 => x"14a9",	130 => x"14d2",	131 => x"14fb",
-- 132 => x"1524",	133 => x"154d",	134 => x"1576",	135 => x"159f",	136 => x"15c8",	137 => x"15f1",
-- 138 => x"161a",	139 => x"1643",	140 => x"166c",	141 => x"1695",	142 => x"16be",	143 => x"16e7",
-- 144 => x"1710",	145 => x"1739",	146 => x"1762",	147 => x"178b",	148 => x"17b4",	149 => x"17dd",
-- 150 => x"1806",	151 => x"182f",	152 => x"1858",	153 => x"1881",	154 => x"18aa",	155 => x"18d3",
-- 156 => x"18fc",	157 => x"1925",	158 => x"194e",	159 => x"1977",	160 => x"19a0",	161 => x"19c9",
-- 162 => x"19f2",	163 => x"1a1b",	164 => x"1a44",	165 => x"1a6d",	166 => x"1a96",	167 => x"1abf",
-- 168 => x"1ae8",	169 => x"1b11",	170 => x"1b3a",	171 => x"1b63",	172 => x"1b8c",	173 => x"1bb5",
-- 174 => x"1bde",	175 => x"1c07",	176 => x"1c30",	177 => x"1c59",	178 => x"1c82",	179 => x"1cab",
-- 180 => x"1cd4",	181 => x"1cfd",	182 => x"1d26",	183 => x"1d4f",	184 => x"1d78",	185 => x"1da1",
-- 186 => x"1dca",	187 => x"1df3",	188 => x"1e1c",	189 => x"1e45",	190 => x"1e6e",	191 => x"1e97",
-- 192 => x"1ec0",	193 => x"1ee9",	194 => x"1f12",	195 => x"1f3b",	196 => x"1f64",	197 => x"1f8d",
-- 198 => x"1fb6",	199 => x"1fdf",	200 => x"2008",	201 => x"2031",	202 => x"205a",	203 => x"2083",
-- 204 => x"20ac",	205 => x"20d5",	206 => x"20fe",	207 => x"2127",	208 => x"2150",	209 => x"2179",
-- 210 => x"21a2",	211 => x"21cb",	212 => x"21f4",	213 => x"221d",	214 => x"2246",	215 => x"226f",
-- 216 => x"2298",	217 => x"22c1",	218 => x"22ea",	219 => x"2313",	220 => x"233c",	221 => x"2365",
-- 222 => x"238e",	223 => x"23b7",	224 => x"23e0",	225 => x"2409",	226 => x"2432",	227 => x"245b",
-- 228 => x"2484",	229 => x"24ad",	230 => x"24d6",	231 => x"24ff",	232 => x"2528",	233 => x"2551",
-- 234 => x"257a",	235 => x"25a3",	236 => x"25cc",	237 => x"25f5",	238 => x"261e",	239 => x"2647",
-- 240 => x"2670",	241 => x"2699",	242 => x"26c2",	243 => x"26eb",	244 => x"2714",	245 => x"273d",
-- 246 => x"2766",	247 => x"278f",	248 => x"27b8",	249 => x"27e1",	250 => x"280a",	251 => x"2833",
-- 252 => x"285c",	253 => x"2885",	254 => x"28ae",	255 => x"28d7");
--
-- -- 7x7
-- constant c_Gaussian_Lut_7_W1: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0001",	2 => x"0002",	3 => x"0003",	4 => x"0004",	5 => x"0005",
-- 6 => x"0006",	7 => x"0007",	8 => x"0008",	9 => x"0009",	10 => x"000a",	11 => x"000b",
-- 12 => x"000c",	13 => x"000d",	14 => x"000e",	15 => x"000f",	16 => x"0010",	17 => x"0011",
-- 18 => x"0012",	19 => x"0013",	20 => x"0014",	21 => x"0015",	22 => x"0016",	23 => x"0017",
-- 24 => x"0018",	25 => x"0019",	26 => x"001a",	27 => x"001b",	28 => x"001c",	29 => x"001d",
-- 30 => x"001e",	31 => x"001f",	32 => x"0020",	33 => x"0021",	34 => x"0022",	35 => x"0023",
-- 36 => x"0024",	37 => x"0025",	38 => x"0026",	39 => x"0027",	40 => x"0028",	41 => x"0029",
-- 42 => x"002a",	43 => x"002b",	44 => x"002c",	45 => x"002d",	46 => x"002e",	47 => x"002f",
-- 48 => x"0030",	49 => x"0031",	50 => x"0032",	51 => x"0033",	52 => x"0034",	53 => x"0035",
-- 54 => x"0036",	55 => x"0037",	56 => x"0038",	57 => x"0039",	58 => x"003a",	59 => x"003b",
-- 60 => x"003c",	61 => x"003d",	62 => x"003e",	63 => x"003f",	64 => x"0040",	65 => x"0041",
-- 66 => x"0042",	67 => x"0043",	68 => x"0044",	69 => x"0045",	70 => x"0046",	71 => x"0047",
-- 72 => x"0048",	73 => x"0049",	74 => x"004a",	75 => x"004b",	76 => x"004c",	77 => x"004d",
-- 78 => x"004e",	79 => x"004f",	80 => x"0050",	81 => x"0051",	82 => x"0052",	83 => x"0053",
-- 84 => x"0054",	85 => x"0055",	86 => x"0056",	87 => x"0057",	88 => x"0058",	89 => x"0059",
-- 90 => x"005a",	91 => x"005b",	92 => x"005c",	93 => x"005d",	94 => x"005e",	95 => x"005f",
-- 96 => x"0060",	97 => x"0061",	98 => x"0062",	99 => x"0063",	100 => x"0064",	101 => x"0065",
-- 102 => x"0066",	103 => x"0067",	104 => x"0068",	105 => x"0069",	106 => x"006a",	107 => x"006b",
-- 108 => x"006c",	109 => x"006d",	110 => x"006e",	111 => x"006f",	112 => x"0070",	113 => x"0071",
-- 114 => x"0072",	115 => x"0073",	116 => x"0074",	117 => x"0075",	118 => x"0076",	119 => x"0077",
-- 120 => x"0078",	121 => x"0079",	122 => x"007a",	123 => x"007b",	124 => x"007c",	125 => x"007d",
-- 126 => x"007e",	127 => x"007f",	128 => x"0080",	129 => x"0081",	130 => x"0082",	131 => x"0083",
-- 132 => x"0084",	133 => x"0085",	134 => x"0086",	135 => x"0087",	136 => x"0088",	137 => x"0089",
-- 138 => x"008a",	139 => x"008b",	140 => x"008c",	141 => x"008d",	142 => x"008e",	143 => x"008f",
-- 144 => x"0090",	145 => x"0091",	146 => x"0092",	147 => x"0093",	148 => x"0094",	149 => x"0095",
-- 150 => x"0096",	151 => x"0097",	152 => x"0098",	153 => x"0099",	154 => x"009a",	155 => x"009b",
-- 156 => x"009c",	157 => x"009d",	158 => x"009e",	159 => x"009f",	160 => x"00a0",	161 => x"00a1",
-- 162 => x"00a2",	163 => x"00a3",	164 => x"00a4",	165 => x"00a5",	166 => x"00a6",	167 => x"00a7",
-- 168 => x"00a8",	169 => x"00a9",	170 => x"00aa",	171 => x"00ab",	172 => x"00ac",	173 => x"00ad",
-- 174 => x"00ae",	175 => x"00af",	176 => x"00b0",	177 => x"00b1",	178 => x"00b2",	179 => x"00b3",
-- 180 => x"00b4",	181 => x"00b5",	182 => x"00b6",	183 => x"00b7",	184 => x"00b8",	185 => x"00b9",
-- 186 => x"00ba",	187 => x"00bb",	188 => x"00bc",	189 => x"00bd",	190 => x"00be",	191 => x"00bf",
-- 192 => x"00c0",	193 => x"00c1",	194 => x"00c2",	195 => x"00c3",	196 => x"00c4",	197 => x"00c5",
-- 198 => x"00c6",	199 => x"00c7",	200 => x"00c8",	201 => x"00c9",	202 => x"00ca",	203 => x"00cb",
-- 204 => x"00cc",	205 => x"00cd",	206 => x"00ce",	207 => x"00cf",	208 => x"00d0",	209 => x"00d1",
-- 210 => x"00d2",	211 => x"00d3",	212 => x"00d4",	213 => x"00d5",	214 => x"00d6",	215 => x"00d7",
-- 216 => x"00d8",	217 => x"00d9",	218 => x"00da",	219 => x"00db",	220 => x"00dc",	221 => x"00dd",
-- 222 => x"00de",	223 => x"00df",	224 => x"00e0",	225 => x"00e1",	226 => x"00e2",	227 => x"00e3",
-- 228 => x"00e4",	229 => x"00e5",	230 => x"00e6",	231 => x"00e7",	232 => x"00e8",	233 => x"00e9",
-- 234 => x"00ea",	235 => x"00eb",	236 => x"00ec",	237 => x"00ed",	238 => x"00ee",	239 => x"00ef",
-- 240 => x"00f0",	241 => x"00f1",	242 => x"00f2",	243 => x"00f3",	244 => x"00f4",	245 => x"00f5",
-- 246 => x"00f6",	247 => x"00f7",	248 => x"00f8",	249 => x"00f9",	250 => x"00fa",	251 => x"00fb",
-- 252 => x"00fc",	253 => x"00fd",	254 => x"00fe",	255 => x"00ff");
--
-- constant c_Gaussian_Lut_7_W2: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0003",	2 => x"0006",	3 => x"0009",	4 => x"000c",	5 => x"000f",
-- 6 => x"0012",	7 => x"0015",	8 => x"0018",	9 => x"001b",	10 => x"001e",	11 => x"0021",
-- 12 => x"0024",	13 => x"0027",	14 => x"002a",	15 => x"002d",	16 => x"0030",	17 => x"0033",
-- 18 => x"0036",	19 => x"0039",	20 => x"003c",	21 => x"003f",	22 => x"0042",	23 => x"0045",
-- 24 => x"0048",	25 => x"004b",	26 => x"004e",	27 => x"0051",	28 => x"0054",	29 => x"0057",
-- 30 => x"005a",	31 => x"005d",	32 => x"0060",	33 => x"0063",	34 => x"0066",	35 => x"0069",
-- 36 => x"006c",	37 => x"006f",	38 => x"0072",	39 => x"0075",	40 => x"0078",	41 => x"007b",
-- 42 => x"007e",	43 => x"0081",	44 => x"0084",	45 => x"0087",	46 => x"008a",	47 => x"008d",
-- 48 => x"0090",	49 => x"0093",	50 => x"0096",	51 => x"0099",	52 => x"009c",	53 => x"009f",
-- 54 => x"00a2",	55 => x"00a5",	56 => x"00a8",	57 => x"00ab",	58 => x"00ae",	59 => x"00b1",
-- 60 => x"00b4",	61 => x"00b7",	62 => x"00ba",	63 => x"00bd",	64 => x"00c0",	65 => x"00c3",
-- 66 => x"00c6",	67 => x"00c9",	68 => x"00cc",	69 => x"00cf",	70 => x"00d2",	71 => x"00d5",
-- 72 => x"00d8",	73 => x"00db",	74 => x"00de",	75 => x"00e1",	76 => x"00e4",	77 => x"00e7",
-- 78 => x"00ea",	79 => x"00ed",	80 => x"00f0",	81 => x"00f3",	82 => x"00f6",	83 => x"00f9",
-- 84 => x"00fc",	85 => x"00ff",	86 => x"0102",	87 => x"0105",	88 => x"0108",	89 => x"010b",
-- 90 => x"010e",	91 => x"0111",	92 => x"0114",	93 => x"0117",	94 => x"011a",	95 => x"011d",
-- 96 => x"0120",	97 => x"0123",	98 => x"0126",	99 => x"0129",	100 => x"012c",	101 => x"012f",
-- 102 => x"0132",	103 => x"0135",	104 => x"0138",	105 => x"013b",	106 => x"013e",	107 => x"0141",
-- 108 => x"0144",	109 => x"0147",	110 => x"014a",	111 => x"014d",	112 => x"0150",	113 => x"0153",
-- 114 => x"0156",	115 => x"0159",	116 => x"015c",	117 => x"015f",	118 => x"0162",	119 => x"0165",
-- 120 => x"0168",	121 => x"016b",	122 => x"016e",	123 => x"0171",	124 => x"0174",	125 => x"0177",
-- 126 => x"017a",	127 => x"017d",	128 => x"0180",	129 => x"0183",	130 => x"0186",	131 => x"0189",
-- 132 => x"018c",	133 => x"018f",	134 => x"0192",	135 => x"0195",	136 => x"0198",	137 => x"019b",
-- 138 => x"019e",	139 => x"01a1",	140 => x"01a4",	141 => x"01a7",	142 => x"01aa",	143 => x"01ad",
-- 144 => x"01b0",	145 => x"01b3",	146 => x"01b6",	147 => x"01b9",	148 => x"01bc",	149 => x"01bf",
-- 150 => x"01c2",	151 => x"01c5",	152 => x"01c8",	153 => x"01cb",	154 => x"01ce",	155 => x"01d1",
-- 156 => x"01d4",	157 => x"01d7",	158 => x"01da",	159 => x"01dd",	160 => x"01e0",	161 => x"01e3",
-- 162 => x"01e6",	163 => x"01e9",	164 => x"01ec",	165 => x"01ef",	166 => x"01f2",	167 => x"01f5",
-- 168 => x"01f8",	169 => x"01fb",	170 => x"01fe",	171 => x"0201",	172 => x"0204",	173 => x"0207",
-- 174 => x"020a",	175 => x"020d",	176 => x"0210",	177 => x"0213",	178 => x"0216",	179 => x"0219",
-- 180 => x"021c",	181 => x"021f",	182 => x"0222",	183 => x"0225",	184 => x"0228",	185 => x"022b",
-- 186 => x"022e",	187 => x"0231",	188 => x"0234",	189 => x"0237",	190 => x"023a",	191 => x"023d",
-- 192 => x"0240",	193 => x"0243",	194 => x"0246",	195 => x"0249",	196 => x"024c",	197 => x"024f",
-- 198 => x"0252",	199 => x"0255",	200 => x"0258",	201 => x"025b",	202 => x"025e",	203 => x"0261",
-- 204 => x"0264",	205 => x"0267",	206 => x"026a",	207 => x"026d",	208 => x"0270",	209 => x"0273",
-- 210 => x"0276",	211 => x"0279",	212 => x"027c",	213 => x"027f",	214 => x"0282",	215 => x"0285",
-- 216 => x"0288",	217 => x"028b",	218 => x"028e",	219 => x"0291",	220 => x"0294",	221 => x"0297",
-- 222 => x"029a",	223 => x"029d",	224 => x"02a0",	225 => x"02a3",	226 => x"02a6",	227 => x"02a9",
-- 228 => x"02ac",	229 => x"02af",	230 => x"02b2",	231 => x"02b5",	232 => x"02b8",	233 => x"02bb",
-- 234 => x"02be",	235 => x"02c1",	236 => x"02c4",	237 => x"02c7",	238 => x"02ca",	239 => x"02cd",
-- 240 => x"02d0",	241 => x"02d3",	242 => x"02d6",	243 => x"02d9",	244 => x"02dc",	245 => x"02df",
-- 246 => x"02e2",	247 => x"02e5",	248 => x"02e8",	249 => x"02eb",	250 => x"02ee",	251 => x"02f1",
-- 252 => x"02f4",	253 => x"02f7",	254 => x"02fa",	255 => x"02fd");
--
-- constant c_Gaussian_Lut_7_W3: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0006",	2 => x"000c",	3 => x"0012",	4 => x"0018",	5 => x"001e",
-- 6 => x"0024",	7 => x"002a",	8 => x"0030",	9 => x"0036",	10 => x"003c",	11 => x"0042",
-- 12 => x"0048",	13 => x"004e",	14 => x"0054",	15 => x"005a",	16 => x"0060",	17 => x"0066",
-- 18 => x"006c",	19 => x"0072",	20 => x"0078",	21 => x"007e",	22 => x"0084",	23 => x"008a",
-- 24 => x"0090",	25 => x"0096",	26 => x"009c",	27 => x"00a2",	28 => x"00a8",	29 => x"00ae",
-- 30 => x"00b4",	31 => x"00ba",	32 => x"00c0",	33 => x"00c6",	34 => x"00cc",	35 => x"00d2",
-- 36 => x"00d8",	37 => x"00de",	38 => x"00e4",	39 => x"00ea",	40 => x"00f0",	41 => x"00f6",
-- 42 => x"00fc",	43 => x"0102",	44 => x"0108",	45 => x"010e",	46 => x"0114",	47 => x"011a",
-- 48 => x"0120",	49 => x"0126",	50 => x"012c",	51 => x"0132",	52 => x"0138",	53 => x"013e",
-- 54 => x"0144",	55 => x"014a",	56 => x"0150",	57 => x"0156",	58 => x"015c",	59 => x"0162",
-- 60 => x"0168",	61 => x"016e",	62 => x"0174",	63 => x"017a",	64 => x"0180",	65 => x"0186",
-- 66 => x"018c",	67 => x"0192",	68 => x"0198",	69 => x"019e",	70 => x"01a4",	71 => x"01aa",
-- 72 => x"01b0",	73 => x"01b6",	74 => x"01bc",	75 => x"01c2",	76 => x"01c8",	77 => x"01ce",
-- 78 => x"01d4",	79 => x"01da",	80 => x"01e0",	81 => x"01e6",	82 => x"01ec",	83 => x"01f2",
-- 84 => x"01f8",	85 => x"01fe",	86 => x"0204",	87 => x"020a",	88 => x"0210",	89 => x"0216",
-- 90 => x"021c",	91 => x"0222",	92 => x"0228",	93 => x"022e",	94 => x"0234",	95 => x"023a",
-- 96 => x"0240",	97 => x"0246",	98 => x"024c",	99 => x"0252",	100 => x"0258",	101 => x"025e",
-- 102 => x"0264",	103 => x"026a",	104 => x"0270",	105 => x"0276",	106 => x"027c",	107 => x"0282",
-- 108 => x"0288",	109 => x"028e",	110 => x"0294",	111 => x"029a",	112 => x"02a0",	113 => x"02a6",
-- 114 => x"02ac",	115 => x"02b2",	116 => x"02b8",	117 => x"02be",	118 => x"02c4",	119 => x"02ca",
-- 120 => x"02d0",	121 => x"02d6",	122 => x"02dc",	123 => x"02e2",	124 => x"02e8",	125 => x"02ee",
-- 126 => x"02f4",	127 => x"02fa",	128 => x"0300",	129 => x"0306",	130 => x"030c",	131 => x"0312",
-- 132 => x"0318",	133 => x"031e",	134 => x"0324",	135 => x"032a",	136 => x"0330",	137 => x"0336",
-- 138 => x"033c",	139 => x"0342",	140 => x"0348",	141 => x"034e",	142 => x"0354",	143 => x"035a",
-- 144 => x"0360",	145 => x"0366",	146 => x"036c",	147 => x"0372",	148 => x"0378",	149 => x"037e",
-- 150 => x"0384",	151 => x"038a",	152 => x"0390",	153 => x"0396",	154 => x"039c",	155 => x"03a2",
-- 156 => x"03a8",	157 => x"03ae",	158 => x"03b4",	159 => x"03ba",	160 => x"03c0",	161 => x"03c6",
-- 162 => x"03cc",	163 => x"03d2",	164 => x"03d8",	165 => x"03de",	166 => x"03e4",	167 => x"03ea",
-- 168 => x"03f0",	169 => x"03f6",	170 => x"03fc",	171 => x"0402",	172 => x"0408",	173 => x"040e",
-- 174 => x"0414",	175 => x"041a",	176 => x"0420",	177 => x"0426",	178 => x"042c",	179 => x"0432",
-- 180 => x"0438",	181 => x"043e",	182 => x"0444",	183 => x"044a",	184 => x"0450",	185 => x"0456",
-- 186 => x"045c",	187 => x"0462",	188 => x"0468",	189 => x"046e",	190 => x"0474",	191 => x"047a",
-- 192 => x"0480",	193 => x"0486",	194 => x"048c",	195 => x"0492",	196 => x"0498",	197 => x"049e",
-- 198 => x"04a4",	199 => x"04aa",	200 => x"04b0",	201 => x"04b6",	202 => x"04bc",	203 => x"04c2",
-- 204 => x"04c8",	205 => x"04ce",	206 => x"04d4",	207 => x"04da",	208 => x"04e0",	209 => x"04e6",
-- 210 => x"04ec",	211 => x"04f2",	212 => x"04f8",	213 => x"04fe",	214 => x"0504",	215 => x"050a",
-- 216 => x"0510",	217 => x"0516",	218 => x"051c",	219 => x"0522",	220 => x"0528",	221 => x"052e",
-- 222 => x"0534",	223 => x"053a",	224 => x"0540",	225 => x"0546",	226 => x"054c",	227 => x"0552",
-- 228 => x"0558",	229 => x"055e",	230 => x"0564",	231 => x"056a",	232 => x"0570",	233 => x"0576",
-- 234 => x"057c",	235 => x"0582",	236 => x"0588",	237 => x"058e",	238 => x"0594",	239 => x"059a",
-- 240 => x"05a0",	241 => x"05a6",	242 => x"05ac",	243 => x"05b2",	244 => x"05b8",	245 => x"05be",
-- 246 => x"05c4",	247 => x"05ca",	248 => x"05d0",	249 => x"05d6",	250 => x"05dc",	251 => x"05e2",
-- 252 => x"05e8",	253 => x"05ee",	254 => x"05f4",	255 => x"05fa");
--
-- constant c_Gaussian_Lut_7_W4: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"000f",	2 => x"001e",	3 => x"002d",	4 => x"003c",	5 => x"004b",
-- 6 => x"005a",	7 => x"0069",	8 => x"0078",	9 => x"0087",	10 => x"0096",	11 => x"00a5",
-- 12 => x"00b4",	13 => x"00c3",	14 => x"00d2",	15 => x"00e1",	16 => x"00f0",	17 => x"00ff",
-- 18 => x"010e",	19 => x"011d",	20 => x"012c",	21 => x"013b",	22 => x"014a",	23 => x"0159",
-- 24 => x"0168",	25 => x"0177",	26 => x"0186",	27 => x"0195",	28 => x"01a4",	29 => x"01b3",
-- 30 => x"01c2",	31 => x"01d1",	32 => x"01e0",	33 => x"01ef",	34 => x"01fe",	35 => x"020d",
-- 36 => x"021c",	37 => x"022b",	38 => x"023a",	39 => x"0249",	40 => x"0258",	41 => x"0267",
-- 42 => x"0276",	43 => x"0285",	44 => x"0294",	45 => x"02a3",	46 => x"02b2",	47 => x"02c1",
-- 48 => x"02d0",	49 => x"02df",	50 => x"02ee",	51 => x"02fd",	52 => x"030c",	53 => x"031b",
-- 54 => x"032a",	55 => x"0339",	56 => x"0348",	57 => x"0357",	58 => x"0366",	59 => x"0375",
-- 60 => x"0384",	61 => x"0393",	62 => x"03a2",	63 => x"03b1",	64 => x"03c0",	65 => x"03cf",
-- 66 => x"03de",	67 => x"03ed",	68 => x"03fc",	69 => x"040b",	70 => x"041a",	71 => x"0429",
-- 72 => x"0438",	73 => x"0447",	74 => x"0456",	75 => x"0465",	76 => x"0474",	77 => x"0483",
-- 78 => x"0492",	79 => x"04a1",	80 => x"04b0",	81 => x"04bf",	82 => x"04ce",	83 => x"04dd",
-- 84 => x"04ec",	85 => x"04fb",	86 => x"050a",	87 => x"0519",	88 => x"0528",	89 => x"0537",
-- 90 => x"0546",	91 => x"0555",	92 => x"0564",	93 => x"0573",	94 => x"0582",	95 => x"0591",
-- 96 => x"05a0",	97 => x"05af",	98 => x"05be",	99 => x"05cd",	100 => x"05dc",	101 => x"05eb",
-- 102 => x"05fa",	103 => x"0609",	104 => x"0618",	105 => x"0627",	106 => x"0636",	107 => x"0645",
-- 108 => x"0654",	109 => x"0663",	110 => x"0672",	111 => x"0681",	112 => x"0690",	113 => x"069f",
-- 114 => x"06ae",	115 => x"06bd",	116 => x"06cc",	117 => x"06db",	118 => x"06ea",	119 => x"06f9",
-- 120 => x"0708",	121 => x"0717",	122 => x"0726",	123 => x"0735",	124 => x"0744",	125 => x"0753",
-- 126 => x"0762",	127 => x"0771",	128 => x"0780",	129 => x"078f",	130 => x"079e",	131 => x"07ad",
-- 132 => x"07bc",	133 => x"07cb",	134 => x"07da",	135 => x"07e9",	136 => x"07f8",	137 => x"0807",
-- 138 => x"0816",	139 => x"0825",	140 => x"0834",	141 => x"0843",	142 => x"0852",	143 => x"0861",
-- 144 => x"0870",	145 => x"087f",	146 => x"088e",	147 => x"089d",	148 => x"08ac",	149 => x"08bb",
-- 150 => x"08ca",	151 => x"08d9",	152 => x"08e8",	153 => x"08f7",	154 => x"0906",	155 => x"0915",
-- 156 => x"0924",	157 => x"0933",	158 => x"0942",	159 => x"0951",	160 => x"0960",	161 => x"096f",
-- 162 => x"097e",	163 => x"098d",	164 => x"099c",	165 => x"09ab",	166 => x"09ba",	167 => x"09c9",
-- 168 => x"09d8",	169 => x"09e7",	170 => x"09f6",	171 => x"0a05",	172 => x"0a14",	173 => x"0a23",
-- 174 => x"0a32",	175 => x"0a41",	176 => x"0a50",	177 => x"0a5f",	178 => x"0a6e",	179 => x"0a7d",
-- 180 => x"0a8c",	181 => x"0a9b",	182 => x"0aaa",	183 => x"0ab9",	184 => x"0ac8",	185 => x"0ad7",
-- 186 => x"0ae6",	187 => x"0af5",	188 => x"0b04",	189 => x"0b13",	190 => x"0b22",	191 => x"0b31",
-- 192 => x"0b40",	193 => x"0b4f",	194 => x"0b5e",	195 => x"0b6d",	196 => x"0b7c",	197 => x"0b8b",
-- 198 => x"0b9a",	199 => x"0ba9",	200 => x"0bb8",	201 => x"0bc7",	202 => x"0bd6",	203 => x"0be5",
-- 204 => x"0bf4",	205 => x"0c03",	206 => x"0c12",	207 => x"0c21",	208 => x"0c30",	209 => x"0c3f",
-- 210 => x"0c4e",	211 => x"0c5d",	212 => x"0c6c",	213 => x"0c7b",	214 => x"0c8a",	215 => x"0c99",
-- 216 => x"0ca8",	217 => x"0cb7",	218 => x"0cc6",	219 => x"0cd5",	220 => x"0ce4",	221 => x"0cf3",
-- 222 => x"0d02",	223 => x"0d11",	224 => x"0d20",	225 => x"0d2f",	226 => x"0d3e",	227 => x"0d4d",
-- 228 => x"0d5c",	229 => x"0d6b",	230 => x"0d7a",	231 => x"0d89",	232 => x"0d98",	233 => x"0da7",
-- 234 => x"0db6",	235 => x"0dc5",	236 => x"0dd4",	237 => x"0de3",	238 => x"0df2",	239 => x"0e01",
-- 240 => x"0e10",	241 => x"0e1f",	242 => x"0e2e",	243 => x"0e3d",	244 => x"0e4c",	245 => x"0e5b",
-- 246 => x"0e6a",	247 => x"0e79",	248 => x"0e88",	249 => x"0e97",	250 => x"0ea6",	251 => x"0eb5",
-- 252 => x"0ec4",	253 => x"0ed3",	254 => x"0ee2",	255 => x"0ef1");
--
-- constant c_Gaussian_Lut_7_W5: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0019",	2 => x"0032",	3 => x"004b",	4 => x"0064",	5 => x"007d",
-- 6 => x"0096",	7 => x"00af",	8 => x"00c8",	9 => x"00e1",	10 => x"00fa",	11 => x"0113",
-- 12 => x"012c",	13 => x"0145",	14 => x"015e",	15 => x"0177",	16 => x"0190",	17 => x"01a9",
-- 18 => x"01c2",	19 => x"01db",	20 => x"01f4",	21 => x"020d",	22 => x"0226",	23 => x"023f",
-- 24 => x"0258",	25 => x"0271",	26 => x"028a",	27 => x"02a3",	28 => x"02bc",	29 => x"02d5",
-- 30 => x"02ee",	31 => x"0307",	32 => x"0320",	33 => x"0339",	34 => x"0352",	35 => x"036b",
-- 36 => x"0384",	37 => x"039d",	38 => x"03b6",	39 => x"03cf",	40 => x"03e8",	41 => x"0401",
-- 42 => x"041a",	43 => x"0433",	44 => x"044c",	45 => x"0465",	46 => x"047e",	47 => x"0497",
-- 48 => x"04b0",	49 => x"04c9",	50 => x"04e2",	51 => x"04fb",	52 => x"0514",	53 => x"052d",
-- 54 => x"0546",	55 => x"055f",	56 => x"0578",	57 => x"0591",	58 => x"05aa",	59 => x"05c3",
-- 60 => x"05dc",	61 => x"05f5",	62 => x"060e",	63 => x"0627",	64 => x"0640",	65 => x"0659",
-- 66 => x"0672",	67 => x"068b",	68 => x"06a4",	69 => x"06bd",	70 => x"06d6",	71 => x"06ef",
-- 72 => x"0708",	73 => x"0721",	74 => x"073a",	75 => x"0753",	76 => x"076c",	77 => x"0785",
-- 78 => x"079e",	79 => x"07b7",	80 => x"07d0",	81 => x"07e9",	82 => x"0802",	83 => x"081b",
-- 84 => x"0834",	85 => x"084d",	86 => x"0866",	87 => x"087f",	88 => x"0898",	89 => x"08b1",
-- 90 => x"08ca",	91 => x"08e3",	92 => x"08fc",	93 => x"0915",	94 => x"092e",	95 => x"0947",
-- 96 => x"0960",	97 => x"0979",	98 => x"0992",	99 => x"09ab",	100 => x"09c4",	101 => x"09dd",
-- 102 => x"09f6",	103 => x"0a0f",	104 => x"0a28",	105 => x"0a41",	106 => x"0a5a",	107 => x"0a73",
-- 108 => x"0a8c",	109 => x"0aa5",	110 => x"0abe",	111 => x"0ad7",	112 => x"0af0",	113 => x"0b09",
-- 114 => x"0b22",	115 => x"0b3b",	116 => x"0b54",	117 => x"0b6d",	118 => x"0b86",	119 => x"0b9f",
-- 120 => x"0bb8",	121 => x"0bd1",	122 => x"0bea",	123 => x"0c03",	124 => x"0c1c",	125 => x"0c35",
-- 126 => x"0c4e",	127 => x"0c67",	128 => x"0c80",	129 => x"0c99",	130 => x"0cb2",	131 => x"0ccb",
-- 132 => x"0ce4",	133 => x"0cfd",	134 => x"0d16",	135 => x"0d2f",	136 => x"0d48",	137 => x"0d61",
-- 138 => x"0d7a",	139 => x"0d93",	140 => x"0dac",	141 => x"0dc5",	142 => x"0dde",	143 => x"0df7",
-- 144 => x"0e10",	145 => x"0e29",	146 => x"0e42",	147 => x"0e5b",	148 => x"0e74",	149 => x"0e8d",
-- 150 => x"0ea6",	151 => x"0ebf",	152 => x"0ed8",	153 => x"0ef1",	154 => x"0f0a",	155 => x"0f23",
-- 156 => x"0f3c",	157 => x"0f55",	158 => x"0f6e",	159 => x"0f87",	160 => x"0fa0",	161 => x"0fb9",
-- 162 => x"0fd2",	163 => x"0feb",	164 => x"1004",	165 => x"101d",	166 => x"1036",	167 => x"104f",
-- 168 => x"1068",	169 => x"1081",	170 => x"109a",	171 => x"10b3",	172 => x"10cc",	173 => x"10e5",
-- 174 => x"10fe",	175 => x"1117",	176 => x"1130",	177 => x"1149",	178 => x"1162",	179 => x"117b",
-- 180 => x"1194",	181 => x"11ad",	182 => x"11c6",	183 => x"11df",	184 => x"11f8",	185 => x"1211",
-- 186 => x"122a",	187 => x"1243",	188 => x"125c",	189 => x"1275",	190 => x"128e",	191 => x"12a7",
-- 192 => x"12c0",	193 => x"12d9",	194 => x"12f2",	195 => x"130b",	196 => x"1324",	197 => x"133d",
-- 198 => x"1356",	199 => x"136f",	200 => x"1388",	201 => x"13a1",	202 => x"13ba",	203 => x"13d3",
-- 204 => x"13ec",	205 => x"1405",	206 => x"141e",	207 => x"1437",	208 => x"1450",	209 => x"1469",
-- 210 => x"1482",	211 => x"149b",	212 => x"14b4",	213 => x"14cd",	214 => x"14e6",	215 => x"14ff",
-- 216 => x"1518",	217 => x"1531",	218 => x"154a",	219 => x"1563",	220 => x"157c",	221 => x"1595",
-- 222 => x"15ae",	223 => x"15c7",	224 => x"15e0",	225 => x"15f9",	226 => x"1612",	227 => x"162b",
-- 228 => x"1644",	229 => x"165d",	230 => x"1676",	231 => x"168f",	232 => x"16a8",	233 => x"16c1",
-- 234 => x"16da",	235 => x"16f3",	236 => x"170c",	237 => x"1725",	238 => x"173e",	239 => x"1757",
-- 240 => x"1770",	241 => x"1789",	242 => x"17a2",	243 => x"17bb",	244 => x"17d4",	245 => x"17ed",
-- 246 => x"1806",	247 => x"181f",	248 => x"1838",	249 => x"1851",	250 => x"186a",	251 => x"1883",
-- 252 => x"189c",	253 => x"18b5",	254 => x"18ce",	255 => x"18e7");
--
-- constant c_Gaussian_Lut_7_W6: fixed_vector(255 downto 0):= (
-- 0 => x"0000",	1 => x"0029",	2 => x"0052",	3 => x"007b",	4 => x"00a4",	5 => x"00cd",
-- 6 => x"00f6",	7 => x"011f",	8 => x"0148",	9 => x"0171",	10 => x"019a",	11 => x"01c3",
-- 12 => x"01ec",	13 => x"0215",	14 => x"023e",	15 => x"0267",	16 => x"0290",	17 => x"02b9",
-- 18 => x"02e2",	19 => x"030b",	20 => x"0334",	21 => x"035d",	22 => x"0386",	23 => x"03af",
-- 24 => x"03d8",	25 => x"0401",	26 => x"042a",	27 => x"0453",	28 => x"047c",	29 => x"04a5",
-- 30 => x"04ce",	31 => x"04f7",	32 => x"0520",	33 => x"0549",	34 => x"0572",	35 => x"059b",
-- 36 => x"05c4",	37 => x"05ed",	38 => x"0616",	39 => x"063f",	40 => x"0668",	41 => x"0691",
-- 42 => x"06ba",	43 => x"06e3",	44 => x"070c",	45 => x"0735",	46 => x"075e",	47 => x"0787",
-- 48 => x"07b0",	49 => x"07d9",	50 => x"0802",	51 => x"082b",	52 => x"0854",	53 => x"087d",
-- 54 => x"08a6",	55 => x"08cf",	56 => x"08f8",	57 => x"0921",	58 => x"094a",	59 => x"0973",
-- 60 => x"099c",	61 => x"09c5",	62 => x"09ee",	63 => x"0a17",	64 => x"0a40",	65 => x"0a69",
-- 66 => x"0a92",	67 => x"0abb",	68 => x"0ae4",	69 => x"0b0d",	70 => x"0b36",	71 => x"0b5f",
-- 72 => x"0b88",	73 => x"0bb1",	74 => x"0bda",	75 => x"0c03",	76 => x"0c2c",	77 => x"0c55",
-- 78 => x"0c7e",	79 => x"0ca7",	80 => x"0cd0",	81 => x"0cf9",	82 => x"0d22",	83 => x"0d4b",
-- 84 => x"0d74",	85 => x"0d9d",	86 => x"0dc6",	87 => x"0def",	88 => x"0e18",	89 => x"0e41",
-- 90 => x"0e6a",	91 => x"0e93",	92 => x"0ebc",	93 => x"0ee5",	94 => x"0f0e",	95 => x"0f37",
-- 96 => x"0f60",	97 => x"0f89",	98 => x"0fb2",	99 => x"0fdb",	100 => x"1004",	101 => x"102d",
-- 102 => x"1056",	103 => x"107f",	104 => x"10a8",	105 => x"10d1",	106 => x"10fa",	107 => x"1123",
-- 108 => x"114c",	109 => x"1175",	110 => x"119e",	111 => x"11c7",	112 => x"11f0",	113 => x"1219",
-- 114 => x"1242",	115 => x"126b",	116 => x"1294",	117 => x"12bd",	118 => x"12e6",	119 => x"130f",
-- 120 => x"1338",	121 => x"1361",	122 => x"138a",	123 => x"13b3",	124 => x"13dc",	125 => x"1405",
-- 126 => x"142e",	127 => x"1457",	128 => x"1480",	129 => x"14a9",	130 => x"14d2",	131 => x"14fb",
-- 132 => x"1524",	133 => x"154d",	134 => x"1576",	135 => x"159f",	136 => x"15c8",	137 => x"15f1",
-- 138 => x"161a",	139 => x"1643",	140 => x"166c",	141 => x"1695",	142 => x"16be",	143 => x"16e7",
-- 144 => x"1710",	145 => x"1739",	146 => x"1762",	147 => x"178b",	148 => x"17b4",	149 => x"17dd",
-- 150 => x"1806",	151 => x"182f",	152 => x"1858",	153 => x"1881",	154 => x"18aa",	155 => x"18d3",
-- 156 => x"18fc",	157 => x"1925",	158 => x"194e",	159 => x"1977",	160 => x"19a0",	161 => x"19c9",
-- 162 => x"19f2",	163 => x"1a1b",	164 => x"1a44",	165 => x"1a6d",	166 => x"1a96",	167 => x"1abf",
-- 168 => x"1ae8",	169 => x"1b11",	170 => x"1b3a",	171 => x"1b63",	172 => x"1b8c",	173 => x"1bb5",
-- 174 => x"1bde",	175 => x"1c07",	176 => x"1c30",	177 => x"1c59",	178 => x"1c82",	179 => x"1cab",
-- 180 => x"1cd4",	181 => x"1cfd",	182 => x"1d26",	183 => x"1d4f",	184 => x"1d78",	185 => x"1da1",
-- 186 => x"1dca",	187 => x"1df3",	188 => x"1e1c",	189 => x"1e45",	190 => x"1e6e",	191 => x"1e97",
-- 192 => x"1ec0",	193 => x"1ee9",	194 => x"1f12",	195 => x"1f3b",	196 => x"1f64",	197 => x"1f8d",
-- 198 => x"1fb6",	199 => x"1fdf",	200 => x"2008",	201 => x"2031",	202 => x"205a",	203 => x"2083",
-- 204 => x"20ac",	205 => x"20d5",	206 => x"20fe",	207 => x"2127",	208 => x"2150",	209 => x"2179",
-- 210 => x"21a2",	211 => x"21cb",	212 => x"21f4",	213 => x"221d",	214 => x"2246",	215 => x"226f",
-- 216 => x"2298",	217 => x"22c1",	218 => x"22ea",	219 => x"2313",	220 => x"233c",	221 => x"2365",
-- 222 => x"238e",	223 => x"23b7",	224 => x"23e0",	225 => x"2409",	226 => x"2432",	227 => x"245b",
-- 228 => x"2484",	229 => x"24ad",	230 => x"24d6",	231 => x"24ff",	232 => x"2528",	233 => x"2551",
-- 234 => x"257a",	235 => x"25a3",	236 => x"25cc",	237 => x"25f5",	238 => x"261e",	239 => x"2647",
-- 240 => x"2670",	241 => x"2699",	242 => x"26c2",	243 => x"26eb",	244 => x"2714",	245 => x"273d",
-- 246 => x"2766",	247 => x"278f",	248 => x"27b8",	249 => x"27e1",	250 => x"280a",	251 => x"2833",
-- 252 => x"285c",	253 => x"2885",	254 => x"28ae",	255 => x"28d7");

-- Separable values (9.8)
constant c_Gaussian_Kernel_3_Hor : fixed_vector(2 downto 0) := (
	0=>"00000000000010011", 1=>"00000000000100000", 2=>"00000000000010011");
constant c_Gaussian_Kernel_3_Ver : fixed_vector(2 downto 0) := (
	0=>"00000000100000000", 1=>"00000000110100110", 2=>"00000000100000000");

	constant c_Gaussian_Kernel_5_Hor : fixed_vector(4 downto 0) := (
		0=>"00000000000001000", 1=>"00000000000100010", 2=>"00000000000111000", 3=>"00000000000100010", 4=>"00000000000001000");
	constant c_Gaussian_Kernel_5_Ver : fixed_vector(4 downto 0) := (
		0=>"00000000000011010", 1=>"00000000001110011", 2=>"00000000010111101", 3=>"00000000001110011", 4=>"00000000000011010");
constant c_Gaussian_Kernel_7_Hor : fixed_vector(6 downto 0) := (
	0=>"00000000000000001", 1=>"00000000000000110", 2=>"00000000000011011", 3=>"00000000000101101", 4=>"00000000000011011", 5=>"00000000000000110", 6=>"00000000000000001");
constant c_Gaussian_Kernel_7_Ver : fixed_vector(6 downto 0) := (
	0=>"00000000000000011", 1=>"00000000000011111", 2=>"00000000010001100", 3=>"00000000011100110", 4=>"00000000010001100", 5=>"00000000000011111", 6=>"00000000000000011");

end Package_Constant;
