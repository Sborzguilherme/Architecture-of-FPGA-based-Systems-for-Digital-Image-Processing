-- megafunction wizard: %ALTFP_CONVERT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_CONVERT 

-- ============================================================
-- File Name: FPU_CONVERT.vhd
-- Megafunction Name(s):
-- 			ALTFP_CONVERT
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_convert CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="INT2FLOAT" ROUNDING="TO_NEAREST" WIDTH_DATA=32 WIDTH_EXP_INPUT=8 WIDTH_EXP_OUTPUT=8 WIDTH_INT=32 WIDTH_MAN_INPUT=23 WIDTH_MAN_OUTPUT=23 WIDTH_RESULT=32 clock dataa result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:24:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:24:SJ cbx_altfp_convert 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_altsyncram 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_abs 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_compare 2018:09:12:13:04:24:SJ cbx_lpm_decode 2018:09:12:13:04:24:SJ cbx_lpm_divide 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_stratixiii 2018:09:12:13:04:24:SJ cbx_stratixv 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" PIPELINE=2 SHIFTDIR="LEFT" SHIFTTYPE="LOGICAL" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = reg 68 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altbarrel_shift_fof IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altbarrel_shift_fof;

 ARCHITECTURE RTL OF FPU_CONVERT_altbarrel_shift_fof IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper2d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec3r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sel_pipec4r1d	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w97w98w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w93w94w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w118w119w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w114w115w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w140w141w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w136w137w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w162w163w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w158w159w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w181w182w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w177w178w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w89w90w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w110w111w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w132w133w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w154w155w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w173w174w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range82w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range104w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range125w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range149w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_dir_w_range168w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range85w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range106w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range128w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range151w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_sel_w_range170w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w118w119w120w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w140w141w142w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w162w163w164w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w181w182w183w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w100w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w121w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w143w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w165w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w184w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w113w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w116w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w135w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w138w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w157w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w160w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w176w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w179w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range91w92w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w95w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_dir_w_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range145w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range167w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range80w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range103w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sbit_w_range123w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_sel_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range185w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_w_smux_w_range144w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w97w98w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w97w(0) AND wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w95w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w93w94w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w93w(0) AND wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range91w92w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w118w119w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w118w(0) AND wire_altbarrel_shift5_w116w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w114w115w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w114w(0) AND wire_altbarrel_shift5_w113w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w140w141w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w140w(0) AND wire_altbarrel_shift5_w138w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w136w137w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w136w(0) AND wire_altbarrel_shift5_w135w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w162w163w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w162w(0) AND wire_altbarrel_shift5_w160w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w158w159w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w158w(0) AND wire_altbarrel_shift5_w157w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w181w182w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w181w(0) AND wire_altbarrel_shift5_w179w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w177w178w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w177w(0) AND wire_altbarrel_shift5_w176w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w89w90w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range85w89w(0) AND wire_altbarrel_shift5_w_sbit_w_range80w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w110w111w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range106w110w(0) AND wire_altbarrel_shift5_w_sbit_w_range103w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w132w133w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range128w132w(0) AND wire_altbarrel_shift5_w_sbit_w_range123w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w154w155w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range151w154w(0) AND wire_altbarrel_shift5_w_sbit_w_range145w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w173w174w(i) <= wire_altbarrel_shift5_w_lg_w_sel_w_range170w173w(0) AND wire_altbarrel_shift5_w_sbit_w_range167w(i);
	END GENERATE loop14;
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w97w(0) <= wire_altbarrel_shift5_w_sel_w_range85w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range82w96w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w93w(0) <= wire_altbarrel_shift5_w_sel_w_range85w(0) AND wire_altbarrel_shift5_w_dir_w_range82w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w118w(0) <= wire_altbarrel_shift5_w_sel_w_range106w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range104w117w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w114w(0) <= wire_altbarrel_shift5_w_sel_w_range106w(0) AND wire_altbarrel_shift5_w_dir_w_range104w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w140w(0) <= wire_altbarrel_shift5_w_sel_w_range128w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range125w139w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w136w(0) <= wire_altbarrel_shift5_w_sel_w_range128w(0) AND wire_altbarrel_shift5_w_dir_w_range125w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w162w(0) <= wire_altbarrel_shift5_w_sel_w_range151w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range149w161w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w158w(0) <= wire_altbarrel_shift5_w_sel_w_range151w(0) AND wire_altbarrel_shift5_w_dir_w_range149w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w181w(0) <= wire_altbarrel_shift5_w_sel_w_range170w(0) AND wire_altbarrel_shift5_w_lg_w_dir_w_range168w180w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w177w(0) <= wire_altbarrel_shift5_w_sel_w_range170w(0) AND wire_altbarrel_shift5_w_dir_w_range168w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range82w96w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range82w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range104w117w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range104w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range125w139w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range125w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range149w161w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range149w(0);
	wire_altbarrel_shift5_w_lg_w_dir_w_range168w180w(0) <= NOT wire_altbarrel_shift5_w_dir_w_range168w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range85w89w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range85w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range106w110w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range106w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range128w132w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range128w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range151w154w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range151w(0);
	wire_altbarrel_shift5_w_lg_w_sel_w_range170w173w(0) <= NOT wire_altbarrel_shift5_w_sel_w_range170w(0);
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w97w98w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w93w94w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w118w119w120w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w118w119w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w114w115w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w140w141w142w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w140w141w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w136w137w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w162w163w164w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w162w163w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w158w159w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w181w182w183w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w181w182w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w177w178w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w100w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range85w89w90w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w121w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range106w118w119w120w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range106w110w111w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w143w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range128w140w141w142w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range128w132w133w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w165w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range151w162w163w164w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range151w154w155w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 31 GENERATE 
		wire_altbarrel_shift5_w184w(i) <= wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_sel_w_range170w181w182w183w(i) OR wire_altbarrel_shift5_w_lg_w_lg_w_sel_w_range170w173w174w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(1) & dir_w(3) & dir_pipe(0) & dir_w(1 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper2d & smux_w(127 DOWNTO 96) & sbit_piper1d & smux_w(63 DOWNTO 0) & data);
	sel_w <= ( sel_pipec4r1d & sel_pipec3r1d & distance(2 DOWNTO 0));
	smux_w <= ( wire_altbarrel_shift5_w184w & wire_altbarrel_shift5_w165w & wire_altbarrel_shift5_w143w & wire_altbarrel_shift5_w121w & wire_altbarrel_shift5_w_lg_w_lg_w_lg_w_lg_w_sel_w_range85w97w98w99w100w);
	wire_altbarrel_shift5_w113w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_altbarrel_shift5_w116w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_altbarrel_shift5_w135w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_altbarrel_shift5_w138w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_altbarrel_shift5_w157w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_altbarrel_shift5_w160w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_altbarrel_shift5_w176w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_altbarrel_shift5_w179w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_altbarrel_shift5_w_w_pad_w_range87w_w_w_sbit_w_range80w_range91w92w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_altbarrel_shift5_w_w_w_sbit_w_range80w_range88w_w_pad_w_range87w95w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_altbarrel_shift5_w_dir_w_range82w(0) <= dir_w(0);
	wire_altbarrel_shift5_w_dir_w_range104w(0) <= dir_w(1);
	wire_altbarrel_shift5_w_dir_w_range125w(0) <= dir_w(2);
	wire_altbarrel_shift5_w_dir_w_range149w(0) <= dir_w(3);
	wire_altbarrel_shift5_w_dir_w_range168w(0) <= dir_w(4);
	wire_altbarrel_shift5_w_sbit_w_range145w <= sbit_w(127 DOWNTO 96);
	wire_altbarrel_shift5_w_sbit_w_range167w <= sbit_w(159 DOWNTO 128);
	wire_altbarrel_shift5_w_sbit_w_range80w <= sbit_w(31 DOWNTO 0);
	wire_altbarrel_shift5_w_sbit_w_range103w <= sbit_w(63 DOWNTO 32);
	wire_altbarrel_shift5_w_sbit_w_range123w <= sbit_w(95 DOWNTO 64);
	wire_altbarrel_shift5_w_sel_w_range85w(0) <= sel_w(0);
	wire_altbarrel_shift5_w_sel_w_range106w(0) <= sel_w(1);
	wire_altbarrel_shift5_w_sel_w_range128w(0) <= sel_w(2);
	wire_altbarrel_shift5_w_sel_w_range151w(0) <= sel_w(3);
	wire_altbarrel_shift5_w_sel_w_range170w(0) <= sel_w(4);
	wire_altbarrel_shift5_w_smux_w_range185w <= smux_w(159 DOWNTO 128);
	wire_altbarrel_shift5_w_smux_w_range144w <= smux_w(95 DOWNTO 64);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe <= ( dir_w(4) & dir_w(2));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_altbarrel_shift5_w_smux_w_range144w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper2d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper2d <= wire_altbarrel_shift5_w_smux_w_range185w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec3r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec3r1d <= distance(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sel_pipec4r1d <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sel_pipec4r1d <= distance(4);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --FPU_CONVERT_altbarrel_shift_fof


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FPU_CONVERT_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --FPU_CONVERT_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FPU_CONVERT_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero221w & wire_altpriority_encoder16_w_lg_w_lg_zero223w224w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  FPU_CONVERT_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	wire_altpriority_encoder16_w_lg_w_lg_zero221w222w(0) <= wire_altpriority_encoder16_w_lg_zero221w(0) AND wire_altpriority_encoder16_q(0);
	wire_altpriority_encoder16_w_lg_zero223w(0) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder16_w_lg_zero221w(0) <= NOT wire_altpriority_encoder16_zero;
	wire_altpriority_encoder16_w_lg_w_lg_zero223w224w(0) <= wire_altpriority_encoder16_w_lg_zero223w(0) OR wire_altpriority_encoder16_w_lg_w_lg_zero221w222w(0);
	altpriority_encoder16 :  FPU_CONVERT_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FPU_CONVERT_altpriority_encoder_be8;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero211w212w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero213w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero213w214w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero211w & wire_altpriority_encoder14_w_lg_w_lg_zero213w214w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  FPU_CONVERT_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop25 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero211w212w(i) <= wire_altpriority_encoder14_w_lg_zero211w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero213w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop26;
	wire_altpriority_encoder14_w_lg_zero211w(0) <= NOT wire_altpriority_encoder14_zero;
	loop27 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero213w214w(i) <= wire_altpriority_encoder14_w_lg_zero213w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero211w212w(i);
	END GENERATE loop27;
	altpriority_encoder14 :  FPU_CONVERT_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END FPU_CONVERT_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero201w202w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero203w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero203w204w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero201w & wire_altpriority_encoder12_w_lg_w_lg_zero203w204w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  FPU_CONVERT_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	loop28 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero201w202w(i) <= wire_altpriority_encoder12_w_lg_zero201w(0) AND wire_altpriority_encoder12_q(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_zero203w(i) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(i);
	END GENERATE loop29;
	wire_altpriority_encoder12_w_lg_zero201w(0) <= NOT wire_altpriority_encoder12_zero;
	loop30 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder12_w_lg_w_lg_zero203w204w(i) <= wire_altpriority_encoder12_w_lg_zero203w(i) OR wire_altpriority_encoder12_w_lg_w_lg_zero201w202w(i);
	END GENERATE loop30;
	altpriority_encoder12 :  FPU_CONVERT_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_rf8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --FPU_CONVERT_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero255w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero257w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero255w & wire_altpriority_encoder22_w_lg_w_lg_zero257w258w);
	altpriority_encoder21 :  FPU_CONVERT_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder21_q
	  );
	wire_altpriority_encoder22_w_lg_w_lg_zero255w256w(0) <= wire_altpriority_encoder22_w_lg_zero255w(0) AND wire_altpriority_encoder22_q(0);
	wire_altpriority_encoder22_w_lg_zero257w(0) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(0);
	wire_altpriority_encoder22_w_lg_zero255w(0) <= NOT wire_altpriority_encoder22_zero;
	wire_altpriority_encoder22_w_lg_w_lg_zero257w258w(0) <= wire_altpriority_encoder22_w_lg_zero257w(0) OR wire_altpriority_encoder22_w_lg_w_lg_zero255w256w(0);
	altpriority_encoder22 :  FPU_CONVERT_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_6v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero246w247w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero248w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero248w249w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero246w & wire_altpriority_encoder20_w_lg_w_lg_zero248w249w);
	altpriority_encoder19 :  FPU_CONVERT_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop31 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero246w247w(i) <= wire_altpriority_encoder20_w_lg_zero246w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_zero248w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop32;
	wire_altpriority_encoder20_w_lg_zero246w(0) <= NOT wire_altpriority_encoder20_zero;
	loop33 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero248w249w(i) <= wire_altpriority_encoder20_w_lg_zero248w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero246w247w(i);
	END GENERATE loop33;
	altpriority_encoder20 :  FPU_CONVERT_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_bv7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altpriority_encoder_r08;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero237w238w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero239w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero239w240w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero237w & wire_altpriority_encoder18_w_lg_w_lg_zero239w240w);
	altpriority_encoder17 :  FPU_CONVERT_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop34 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero237w238w(i) <= wire_altpriority_encoder18_w_lg_zero237w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_zero239w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop35;
	wire_altpriority_encoder18_w_lg_zero237w(0) <= NOT wire_altpriority_encoder18_zero;
	loop36 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero239w240w(i) <= wire_altpriority_encoder18_w_lg_zero239w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero237w238w(i);
	END GENERATE loop36;
	altpriority_encoder18 :  FPU_CONVERT_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_r08

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF FPU_CONVERT_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero192w193w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero194w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero194w195w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 COMPONENT  FPU_CONVERT_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero192w & wire_altpriority_encoder10_w_lg_w_lg_zero194w195w);
	loop37 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero192w193w(i) <= wire_altpriority_encoder10_w_lg_zero192w(0) AND wire_altpriority_encoder10_q(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_zero194w(i) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(i);
	END GENERATE loop38;
	wire_altpriority_encoder10_w_lg_zero192w(0) <= NOT wire_altpriority_encoder10_zero;
	loop39 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder10_w_lg_w_lg_zero194w195w(i) <= wire_altpriority_encoder10_w_lg_zero194w(i) OR wire_altpriority_encoder10_w_lg_w_lg_zero192w193w(i);
	END GENERATE loop39;
	altpriority_encoder10 :  FPU_CONVERT_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  FPU_CONVERT_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --FPU_CONVERT_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 5 lpm_compare 1 reg 247 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  FPU_CONVERT_altfp_convert_7qm IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END FPU_CONVERT_altfp_convert_7qm;

 ARCHITECTURE RTL OF FPU_CONVERT_altfp_convert_7qm IS

	 SIGNAL  wire_altbarrel_shift5_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altbarrel_shift5_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 add_1_adder1_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q58w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_1_adder1_cout_reg_w_lg_q60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_1_adder1_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_cout_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_adder2_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 add_1_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_1_reg_w_lg_w_lg_q67w68w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q66w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_1_reg_w_lg_q67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exponent_bus_pre_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponent_bus_pre_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mag_int_a_reg2	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissa_pre_round_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissa_pre_round_reg_w_q_range59w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL	 priority_encoder_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_int_a_reg5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub6_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_cout	:	STD_LOGIC;
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_w_lg_alb21w22w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb20w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_cmpr4_w_lg_alb21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cmpr4_alb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_w52w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mantissa_overflow71w72w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_max_neg_value_selector17w18w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sign_int_a5w6w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow70w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector16w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a4w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mantissa_overflow71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_max_neg_value_selector17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sign_int_a5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range34w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range38w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range41w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range44w46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_or_w_range47w49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_adder1_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder2_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  add_1_adder_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  const_bias_value_add_width_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exceptions_value :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_bus_pre :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_output_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_rounded :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exponent_zero_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  int_a_2s :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  invert_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  leading_zeroes :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mag_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  mantissa_bus :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  mantissa_overflow :	STD_LOGIC;
	 SIGNAL  mantissa_post_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_pre_round :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mantissa_rounded :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  max_neg_value_selector :	STD_LOGIC;
	 SIGNAL  max_neg_value_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  minus_leading_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  prio_mag_int_a :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  shifted_mag_int_a :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  sign_bus :	STD_LOGIC;
	 SIGNAL  sign_int_a :	STD_LOGIC;
	 SIGNAL  sticky_bit_bus :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_or_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  zero_padding_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_bus_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_or_w_range47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  FPU_CONVERT_altbarrel_shift_fof
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  FPU_CONVERT_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w(0) <= wire_w_lg_w_lg_guard_bit_w52w53w(0) AND sticky_bit_w;
	wire_w_lg_w_lg_guard_bit_w52w53w(0) <= wire_w_lg_guard_bit_w52w(0) AND round_bit_w;
	loop40 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_mantissa_overflow71w72w(i) <= wire_w_lg_mantissa_overflow71w(0) AND exponent_bus_pre_reg(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_max_neg_value_selector17w18w(i) <= wire_w_lg_max_neg_value_selector17w(0) AND exponent_zero_w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_sign_int_a5w6w(i) <= wire_w_lg_sign_int_a5w(0) AND int_a(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_mantissa_overflow70w(i) <= mantissa_overflow AND wire_add_sub8_result(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_max_neg_value_selector16w(i) <= max_neg_value_selector AND max_neg_value_w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_sign_int_a4w(i) <= sign_int_a AND int_a_2s(i);
	END GENERATE loop45;
	wire_w_lg_guard_bit_w52w(0) <= NOT guard_bit_w;
	wire_w_lg_mantissa_overflow71w(0) <= NOT mantissa_overflow;
	wire_w_lg_max_neg_value_selector17w(0) <= NOT max_neg_value_selector;
	wire_w_lg_sign_int_a5w(0) <= NOT sign_int_a;
	wire_w_lg_w_sticky_bit_or_w_range34w37w(0) <= wire_w_sticky_bit_or_w_range34w(0) OR wire_w_sticky_bit_bus_range36w(0);
	wire_w_lg_w_sticky_bit_or_w_range38w40w(0) <= wire_w_sticky_bit_or_w_range38w(0) OR wire_w_sticky_bit_bus_range39w(0);
	wire_w_lg_w_sticky_bit_or_w_range41w43w(0) <= wire_w_sticky_bit_or_w_range41w(0) OR wire_w_sticky_bit_bus_range42w(0);
	wire_w_lg_w_sticky_bit_or_w_range44w46w(0) <= wire_w_sticky_bit_or_w_range44w(0) OR wire_w_sticky_bit_bus_range45w(0);
	wire_w_lg_w_sticky_bit_or_w_range47w49w(0) <= wire_w_sticky_bit_or_w_range47w(0) OR wire_w_sticky_bit_bus_range48w(0);
	aclr <= '0';
	add_1_adder1_w <= add_1_adder1_reg;
	add_1_adder2_w <= (wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w OR wire_add_1_adder1_cout_reg_w_lg_q58w);
	add_1_adder_w <= ( add_1_adder2_w & add_1_adder1_w);
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_w52w53w54w(0) OR (guard_bit_w AND round_bit_w));
	bias_value_w <= "01111111";
	clk_en <= '1';
	const_bias_value_add_width_int_w <= "10011101";
	exceptions_value <= (wire_w_lg_w_lg_max_neg_value_selector17w18w OR wire_w_lg_max_neg_value_selector16w);
	exponent_bus <= exponent_rounded;
	exponent_bus_pre <= (wire_cmpr4_w_lg_w_lg_alb21w22w OR wire_cmpr4_w_lg_alb20w);
	exponent_output_w <= wire_add_sub3_result;
	exponent_rounded <= (wire_w_lg_w_lg_mantissa_overflow71w72w OR wire_w_lg_mantissa_overflow70w);
	exponent_zero_w <= (OTHERS => '0');
	guard_bit_w <= shifted_mag_int_a(7);
	int_a <= dataa(30 DOWNTO 0);
	int_a_2s <= wire_add_sub1_result;
	invert_int_a <= (NOT int_a);
	leading_zeroes <= (NOT priority_encoder_reg);
	mag_int_a <= (wire_w_lg_w_lg_sign_int_a5w6w OR wire_w_lg_sign_int_a4w);
	mantissa_bus <= mantissa_rounded(22 DOWNTO 0);
	mantissa_overflow <= ((add_1_reg AND add_1_adder1_cout_reg) AND add_1_adder2_cout_reg);
	mantissa_post_round <= add_1_adder_w;
	mantissa_pre_round <= shifted_mag_int_a(30 DOWNTO 7);
	mantissa_rounded <= (wire_add_1_reg_w_lg_w_lg_q67w68w OR wire_add_1_reg_w_lg_q66w);
	max_neg_value_selector <= (wire_cmpr4_alb AND sign_int_a_reg2);
	max_neg_value_w <= "10011110";
	minus_leading_zero <= ( zero_padding_w & leading_zeroes);
	prio_mag_int_a <= ( mag_int_a_reg & "1");
	result <= result_reg;
	result_w <= ( sign_bus & exponent_bus & mantissa_bus);
	round_bit_w <= shifted_mag_int_a(6);
	shifted_mag_int_a <= wire_altbarrel_shift5_result(30 DOWNTO 0);
	sign_bus <= sign_int_a_reg5;
	sign_int_a <= dataa(31);
	sticky_bit_bus <= shifted_mag_int_a(5 DOWNTO 0);
	sticky_bit_or_w <= ( wire_w_lg_w_sticky_bit_or_w_range47w49w & wire_w_lg_w_sticky_bit_or_w_range44w46w & wire_w_lg_w_sticky_bit_or_w_range41w43w & wire_w_lg_w_sticky_bit_or_w_range38w40w & wire_w_lg_w_sticky_bit_or_w_range34w37w & sticky_bit_bus(0));
	sticky_bit_w <= sticky_bit_or_w(5);
	zero_padding_w <= (OTHERS => '0');
	wire_w_sticky_bit_bus_range36w(0) <= sticky_bit_bus(1);
	wire_w_sticky_bit_bus_range39w(0) <= sticky_bit_bus(2);
	wire_w_sticky_bit_bus_range42w(0) <= sticky_bit_bus(3);
	wire_w_sticky_bit_bus_range45w(0) <= sticky_bit_bus(4);
	wire_w_sticky_bit_bus_range48w(0) <= sticky_bit_bus(5);
	wire_w_sticky_bit_or_w_range34w(0) <= sticky_bit_or_w(0);
	wire_w_sticky_bit_or_w_range38w(0) <= sticky_bit_or_w(1);
	wire_w_sticky_bit_or_w_range41w(0) <= sticky_bit_or_w(2);
	wire_w_sticky_bit_or_w_range44w(0) <= sticky_bit_or_w(3);
	wire_w_sticky_bit_or_w_range47w(0) <= sticky_bit_or_w(4);
	wire_altbarrel_shift5_data <= ( "0" & mag_int_a_reg2);
	altbarrel_shift5 :  FPU_CONVERT_altbarrel_shift_fof
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_altbarrel_shift5_data,
		distance => leading_zeroes,
		result => wire_altbarrel_shift5_result
	  );
	altpriority_encoder2 :  FPU_CONVERT_altpriority_encoder_qb6
	  PORT MAP ( 
		data => prio_mag_int_a,
		q => wire_altpriority_encoder2_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_cout_reg <= wire_add_sub6_cout;
			END IF;
		END IF;
	END PROCESS;
	loop46 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_w_lg_q60w61w(i) <= wire_add_1_adder1_cout_reg_w_lg_q60w(0) AND wire_mantissa_pre_round_reg_w_q_range59w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 11 GENERATE 
		wire_add_1_adder1_cout_reg_w_lg_q58w(i) <= add_1_adder1_cout_reg AND add_1_adder2_reg(i);
	END GENERATE loop47;
	wire_add_1_adder1_cout_reg_w_lg_q60w(0) <= NOT add_1_adder1_cout_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder1_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder1_reg <= wire_add_sub6_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_cout_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_cout_reg <= wire_add_sub7_cout;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_adder2_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_adder2_reg <= wire_add_sub7_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN add_1_reg <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN add_1_reg <= add_1_w;
			END IF;
		END IF;
	END PROCESS;
	loop48 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_w_lg_q67w68w(i) <= wire_add_1_reg_w_lg_q67w(0) AND mantissa_pre_round_reg(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 23 GENERATE 
		wire_add_1_reg_w_lg_q66w(i) <= add_1_reg AND mantissa_post_round(i);
	END GENERATE loop49;
	wire_add_1_reg_w_lg_q67w(0) <= NOT add_1_reg;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg <= exponent_bus_pre_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg2 <= exponent_bus_pre_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponent_bus_pre_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponent_bus_pre_reg3 <= exponent_bus_pre;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg <= mag_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mag_int_a_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mag_int_a_reg2 <= mag_int_a_reg;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissa_pre_round_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissa_pre_round_reg <= mantissa_pre_round;
			END IF;
		END IF;
	END PROCESS;
	wire_mantissa_pre_round_reg_w_q_range59w <= mantissa_pre_round_reg(23 DOWNTO 12);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN priority_encoder_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN priority_encoder_reg <= wire_altpriority_encoder2_q;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_reg <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_reg <= result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg1 <= sign_int_a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg2 <= sign_int_a_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg3 <= sign_int_a_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg4 <= sign_int_a_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_int_a_reg5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_int_a_reg5 <= sign_int_a_reg4;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_datab <= "0000000000000000000000000000001";
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 31,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => invert_int_a,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => const_bias_value_add_width_int_w,
		datab => minus_leading_zero,
		result => wire_add_sub3_result
	  );
	wire_add_sub6_datab <= "000000000001";
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub6_cout,
		dataa => mantissa_pre_round(11 DOWNTO 0),
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	wire_add_sub7_datab <= "000000000001";
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 12,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		cout => wire_add_sub7_cout,
		dataa => mantissa_pre_round(23 DOWNTO 12),
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	wire_add_sub8_datab <= "00000001";
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_WIDTH => 8,
		lpm_hint => "ONE_INPUT_IS_CONSTANT=YES"
	  )
	  PORT MAP ( 
		dataa => exponent_bus_pre_reg,
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	loop50 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_w_lg_alb21w22w(i) <= wire_cmpr4_w_lg_alb21w(0) AND exponent_output_w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 7 GENERATE 
		wire_cmpr4_w_lg_alb20w(i) <= wire_cmpr4_alb AND exceptions_value(i);
	END GENERATE loop51;
	wire_cmpr4_w_lg_alb21w(0) <= NOT wire_cmpr4_alb;
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		alb => wire_cmpr4_alb,
		dataa => exponent_output_w,
		datab => bias_value_w
	  );

 END RTL; --FPU_CONVERT_altfp_convert_7qm
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FPU_CONVERT IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END FPU_CONVERT;


ARCHITECTURE RTL OF fpu_convert IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT FPU_CONVERT_altfp_convert_7qm
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	FPU_CONVERT_altfp_convert_7qm_component : FPU_CONVERT_altfp_convert_7qm
	PORT MAP (
		clock => clock,
		dataa => dataa,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_convert"
-- Retrieval info: CONSTANT: OPERATION STRING "INT2FLOAT"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_DATA NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_EXP_INPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_EXP_OUTPUT NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_INT NUMERIC "32"
-- Retrieval info: CONSTANT: WIDTH_MAN_INPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_MAN_OUTPUT NUMERIC "23"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "32"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT_inst.vhd FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL FPU_CONVERT.cmp FALSE TRUE
-- Retrieval info: LIB_FILE: lpm
